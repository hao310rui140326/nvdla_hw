// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_CSC_pra_cell.v

module CSC_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/CSC_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module CSC_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/CSC_mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module CSC_mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_shift_l_beh_v2.v 
module CSC_mgc_shift_l(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   assign z = signd_a ? fshl_u(a,s,a[width_a-1]) : fshl_u(a,s,1'b0);

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_shift_bl_beh_v2.v 
module CSC_mgc_shift_bl(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   assign z = signd_a ? fshl_s(a,s,a[width_a-1]) : fshl_s(a,s,1'b0);

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_shift_r_beh_v2.v 
module CSC_mgc_shift_r(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   assign z = signd_a ? fshr_u(a,s,a[width_a-1]) : fshr_u(a,s,1'b0);

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-081
//  Generated date: Wed May 17 17:57:36 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    CSC_leading_sign_10_0
// ------------------------------------------------------------------


module CSC_leading_sign_10_0 (
  mantissa, rtn
);
  input [9:0] mantissa;
  output [3:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_3;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc;

  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl;
  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl;
  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[7:6]!=2'b00));
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[9:8]!=2'b00));
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_2 = IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[3:2]==2'b00)
      & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_3 = c_h_1_2 & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc = (mantissa[1:0]==2'b00)
      & c_h_1_3;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl = c_h_1_2 & (~ IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3);
  assign IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl
      = (IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 & (IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1
      | (~ IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2)) & (~ c_h_1_3))
      | IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl
      = ~((mantissa[9]) | (~((mantissa[8:7]!=2'b01))) | (((mantissa[5]) | (~((mantissa[4:3]!=2'b01))))
      & c_h_1_2) | ((mantissa[1]) & c_h_1_3) | IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc);
  assign rtn = {c_h_1_3 , (IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl) , (IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl)
      , (IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl)};
endmodule




//------> ../td_ccore_solutions/leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-147
//  Generated date: Fri Feb 17 16:45:25 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    CSC_leading_sign_23_0
// ------------------------------------------------------------------


module CSC_leading_sign_23_0 (
  mantissa, rtn
);
  input [22:0] mantissa;
  output [4:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_10;

  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[20:19]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[18:17]!=2'b00));
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[16:15]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[12:11]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[10:9]!=2'b00));
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[8:7]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[4:3]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4);
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = c_h_1_2 & (c_h_1_5 | (~
      IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3)) & (c_h_1_9 | (~ c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2)))) & c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl
      = ((~((mantissa[22]) | (~((mantissa[21:20]!=2'b01))))) & (~(((mantissa[18])
      | (~((mantissa[17:16]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[14]) | (~((mantissa[13:12]!=2'b01)))))
      & (~(((mantissa[10]) | (~((mantissa[9:8]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[6]) | (~((mantissa[5:4]!=2'b01))))) & (~((~((mantissa[2:1]==2'b01)))
      & c_h_1_9)))) & c_h_1_10))) | ((~ (mantissa[0])) & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      & c_h_1_9 & c_h_1_10);
  assign rtn = {c_h_1_10 , (IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl)
      , (IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl)};
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-179
//  Generated date: Fri Jun 16 23:44:23 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    CSC_chn_data_out_rsci_unreg
// ------------------------------------------------------------------


module CSC_chn_data_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CSC_chn_data_in_rsci_unreg
// ------------------------------------------------------------------


module CSC_chn_data_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for NV_NVDLA_CSC_pra_cell_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : NV_NVDLA_CSC_pra_cell_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_staller
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_data_in_rsci_wen_comp, core_wten,
      chn_data_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_data_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_data_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_data_in_rsci_wen_comp & chn_data_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_dp
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_data_out_rsci_oswt, chn_data_out_rsci_bawt,
      chn_data_out_rsci_wen_comp, chn_data_out_rsci_biwt, chn_data_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_data_out_rsci_oswt;
  output chn_data_out_rsci_bawt;
  output chn_data_out_rsci_wen_comp;
  input chn_data_out_rsci_biwt;
  input chn_data_out_rsci_bdwt;


  // Interconnect Declarations
  reg chn_data_out_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_data_out_rsci_bawt = chn_data_out_rsci_biwt | chn_data_out_rsci_bcwt;
  assign chn_data_out_rsci_wen_comp = (~ chn_data_out_rsci_oswt) | chn_data_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_data_out_rsci_bcwt <= ~((~(chn_data_out_rsci_bcwt | chn_data_out_rsci_biwt))
          | chn_data_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_ctrl
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_data_out_rsci_oswt, core_wen, core_wten, chn_data_out_rsci_iswt0,
      chn_data_out_rsci_ld_core_psct, chn_data_out_rsci_biwt, chn_data_out_rsci_bdwt,
      chn_data_out_rsci_ld_core_sct, chn_data_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_data_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_data_out_rsci_iswt0;
  input chn_data_out_rsci_ld_core_psct;
  output chn_data_out_rsci_biwt;
  output chn_data_out_rsci_bdwt;
  output chn_data_out_rsci_ld_core_sct;
  input chn_data_out_rsci_vd;


  // Interconnect Declarations
  wire chn_data_out_rsci_ogwt;
  wire chn_data_out_rsci_pdswt0;
  reg chn_data_out_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_data_out_rsci_pdswt0 = (~ core_wten) & chn_data_out_rsci_iswt0;
  assign chn_data_out_rsci_biwt = chn_data_out_rsci_ogwt & chn_data_out_rsci_vd;
  assign chn_data_out_rsci_ogwt = chn_data_out_rsci_pdswt0 | chn_data_out_rsci_icwt;
  assign chn_data_out_rsci_bdwt = chn_data_out_rsci_oswt & core_wen;
  assign chn_data_out_rsci_ld_core_sct = chn_data_out_rsci_ld_core_psct & chn_data_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_data_out_rsci_icwt <= ~((~(chn_data_out_rsci_icwt | chn_data_out_rsci_pdswt0))
          | chn_data_out_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_dp
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsci_oswt, chn_data_in_rsci_bawt,
      chn_data_in_rsci_wen_comp, chn_data_in_rsci_d_mxwt, chn_data_in_rsci_biwt,
      chn_data_in_rsci_bdwt, chn_data_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_data_in_rsci_oswt;
  output chn_data_in_rsci_bawt;
  output chn_data_in_rsci_wen_comp;
  output [255:0] chn_data_in_rsci_d_mxwt;
  input chn_data_in_rsci_biwt;
  input chn_data_in_rsci_bdwt;
  input [255:0] chn_data_in_rsci_d;


  // Interconnect Declarations
  reg chn_data_in_rsci_bcwt;
  reg [255:0] chn_data_in_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_data_in_rsci_bawt = chn_data_in_rsci_biwt | chn_data_in_rsci_bcwt;
  assign chn_data_in_rsci_wen_comp = (~ chn_data_in_rsci_oswt) | chn_data_in_rsci_bawt;
  assign chn_data_in_rsci_d_mxwt = MUX_v_256_2_2(chn_data_in_rsci_d, chn_data_in_rsci_d_bfwt,
      chn_data_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_in_rsci_bcwt <= 1'b0;
      chn_data_in_rsci_d_bfwt <= 256'b0;
    end
    else begin
      chn_data_in_rsci_bcwt <= ~((~(chn_data_in_rsci_bcwt | chn_data_in_rsci_biwt))
          | chn_data_in_rsci_bdwt);
      chn_data_in_rsci_d_bfwt <= chn_data_in_rsci_d_mxwt;
    end
  end

  function [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_ctrl
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsci_oswt, core_wen, chn_data_in_rsci_iswt0,
      chn_data_in_rsci_ld_core_psct, core_wten, chn_data_in_rsci_biwt, chn_data_in_rsci_bdwt,
      chn_data_in_rsci_ld_core_sct, chn_data_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_data_in_rsci_oswt;
  input core_wen;
  input chn_data_in_rsci_iswt0;
  input chn_data_in_rsci_ld_core_psct;
  input core_wten;
  output chn_data_in_rsci_biwt;
  output chn_data_in_rsci_bdwt;
  output chn_data_in_rsci_ld_core_sct;
  input chn_data_in_rsci_vd;


  // Interconnect Declarations
  wire chn_data_in_rsci_ogwt;
  wire chn_data_in_rsci_pdswt0;
  reg chn_data_in_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_data_in_rsci_pdswt0 = (~ core_wten) & chn_data_in_rsci_iswt0;
  assign chn_data_in_rsci_biwt = chn_data_in_rsci_ogwt & chn_data_in_rsci_vd;
  assign chn_data_in_rsci_ogwt = chn_data_in_rsci_pdswt0 | chn_data_in_rsci_icwt;
  assign chn_data_in_rsci_bdwt = chn_data_in_rsci_oswt & core_wen;
  assign chn_data_in_rsci_ld_core_sct = chn_data_in_rsci_ld_core_psct & chn_data_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_data_in_rsci_icwt <= ~((~(chn_data_in_rsci_icwt | chn_data_in_rsci_pdswt0))
          | chn_data_in_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_data_out_rsc_z, chn_data_out_rsc_vz, chn_data_out_rsc_lz,
      chn_data_out_rsci_oswt, core_wen, core_wten, chn_data_out_rsci_iswt0, chn_data_out_rsci_bawt,
      chn_data_out_rsci_wen_comp, chn_data_out_rsci_ld_core_psct, chn_data_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [255:0] chn_data_out_rsc_z;
  input chn_data_out_rsc_vz;
  output chn_data_out_rsc_lz;
  input chn_data_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_data_out_rsci_iswt0;
  output chn_data_out_rsci_bawt;
  output chn_data_out_rsci_wen_comp;
  input chn_data_out_rsci_ld_core_psct;
  input [255:0] chn_data_out_rsci_d;


  // Interconnect Declarations
  wire chn_data_out_rsci_biwt;
  wire chn_data_out_rsci_bdwt;
  wire chn_data_out_rsci_ld_core_sct;
  wire chn_data_out_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  CSC_mgc_out_stdreg_wait_v1 #(.rscid(32'sd4),
  .width(32'sd256)) chn_data_out_rsci (
      .ld(chn_data_out_rsci_ld_core_sct),
      .vd(chn_data_out_rsci_vd),
      .d(chn_data_out_rsci_d),
      .lz(chn_data_out_rsc_lz),
      .vz(chn_data_out_rsc_vz),
      .z(chn_data_out_rsc_z)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_ctrl NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_out_rsci_oswt(chn_data_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_data_out_rsci_iswt0(chn_data_out_rsci_iswt0),
      .chn_data_out_rsci_ld_core_psct(chn_data_out_rsci_ld_core_psct),
      .chn_data_out_rsci_biwt(chn_data_out_rsci_biwt),
      .chn_data_out_rsci_bdwt(chn_data_out_rsci_bdwt),
      .chn_data_out_rsci_ld_core_sct(chn_data_out_rsci_ld_core_sct),
      .chn_data_out_rsci_vd(chn_data_out_rsci_vd)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_dp NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_chn_data_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_out_rsci_oswt(chn_data_out_rsci_oswt),
      .chn_data_out_rsci_bawt(chn_data_out_rsci_bawt),
      .chn_data_out_rsci_wen_comp(chn_data_out_rsci_wen_comp),
      .chn_data_out_rsci_biwt(chn_data_out_rsci_biwt),
      .chn_data_out_rsci_bdwt(chn_data_out_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsc_z, chn_data_in_rsc_vz, chn_data_in_rsc_lz,
      chn_data_in_rsci_oswt, core_wen, chn_data_in_rsci_iswt0, chn_data_in_rsci_bawt,
      chn_data_in_rsci_wen_comp, chn_data_in_rsci_ld_core_psct, chn_data_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [255:0] chn_data_in_rsc_z;
  input chn_data_in_rsc_vz;
  output chn_data_in_rsc_lz;
  input chn_data_in_rsci_oswt;
  input core_wen;
  input chn_data_in_rsci_iswt0;
  output chn_data_in_rsci_bawt;
  output chn_data_in_rsci_wen_comp;
  input chn_data_in_rsci_ld_core_psct;
  output [255:0] chn_data_in_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_data_in_rsci_biwt;
  wire chn_data_in_rsci_bdwt;
  wire chn_data_in_rsci_ld_core_sct;
  wire chn_data_in_rsci_vd;
  wire [255:0] chn_data_in_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  CSC_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd256)) chn_data_in_rsci (
      .ld(chn_data_in_rsci_ld_core_sct),
      .vd(chn_data_in_rsci_vd),
      .d(chn_data_in_rsci_d),
      .lz(chn_data_in_rsc_lz),
      .vz(chn_data_in_rsc_vz),
      .z(chn_data_in_rsc_z)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_ctrl NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_in_rsci_oswt(chn_data_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_data_in_rsci_iswt0(chn_data_in_rsci_iswt0),
      .chn_data_in_rsci_ld_core_psct(chn_data_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_data_in_rsci_biwt(chn_data_in_rsci_biwt),
      .chn_data_in_rsci_bdwt(chn_data_in_rsci_bdwt),
      .chn_data_in_rsci_ld_core_sct(chn_data_in_rsci_ld_core_sct),
      .chn_data_in_rsci_vd(chn_data_in_rsci_vd)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_dp NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_chn_data_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_in_rsci_oswt(chn_data_in_rsci_oswt),
      .chn_data_in_rsci_bawt(chn_data_in_rsci_bawt),
      .chn_data_in_rsci_wen_comp(chn_data_in_rsci_wen_comp),
      .chn_data_in_rsci_d_mxwt(chn_data_in_rsci_d_mxwt),
      .chn_data_in_rsci_biwt(chn_data_in_rsci_biwt),
      .chn_data_in_rsci_bdwt(chn_data_in_rsci_bdwt),
      .chn_data_in_rsci_d(chn_data_in_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell_core
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell_core (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsc_z, chn_data_in_rsc_vz, chn_data_in_rsc_lz,
      cfg_precision, cfg_truncate_rsc_z, chn_data_out_rsc_z, chn_data_out_rsc_vz,
      chn_data_out_rsc_lz, chn_data_in_rsci_oswt, chn_data_in_rsci_oswt_unreg, chn_data_out_rsci_oswt,
      chn_data_out_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [255:0] chn_data_in_rsc_z;
  input chn_data_in_rsc_vz;
  output chn_data_in_rsc_lz;
  input [1:0] cfg_precision;
  input [1:0] cfg_truncate_rsc_z;
  output [255:0] chn_data_out_rsc_z;
  input chn_data_out_rsc_vz;
  output chn_data_out_rsc_lz;
  input chn_data_in_rsci_oswt;
  output chn_data_in_rsci_oswt_unreg;
  input chn_data_out_rsci_oswt;
  output chn_data_out_rsci_oswt_unreg;


  // Interconnect Declarations
  wire core_wen;
  reg chn_data_in_rsci_iswt0;
  wire chn_data_in_rsci_bawt;
  wire chn_data_in_rsci_wen_comp;
  reg chn_data_in_rsci_ld_core_psct;
  wire [255:0] chn_data_in_rsci_d_mxwt;
  wire core_wten;
  wire [1:0] cfg_truncate_rsci_d;
  reg chn_data_out_rsci_iswt0;
  wire chn_data_out_rsci_bawt;
  wire chn_data_out_rsci_wen_comp;
  reg chn_data_out_rsci_d_255;
  reg chn_data_out_rsci_d_254;
  reg [3:0] chn_data_out_rsci_d_253_250;
  reg [2:0] chn_data_out_rsci_d_249_247;
  reg [5:0] chn_data_out_rsci_d_246_241;
  reg chn_data_out_rsci_d_240;
  reg chn_data_out_rsci_d_239;
  reg chn_data_out_rsci_d_238;
  reg [3:0] chn_data_out_rsci_d_237_234;
  reg [2:0] chn_data_out_rsci_d_233_231;
  reg [5:0] chn_data_out_rsci_d_230_225;
  reg chn_data_out_rsci_d_224;
  reg chn_data_out_rsci_d_223;
  reg chn_data_out_rsci_d_222;
  reg [3:0] chn_data_out_rsci_d_221_218;
  reg [2:0] chn_data_out_rsci_d_217_215;
  reg [5:0] chn_data_out_rsci_d_214_209;
  reg chn_data_out_rsci_d_208;
  reg chn_data_out_rsci_d_207;
  reg chn_data_out_rsci_d_206;
  reg [3:0] chn_data_out_rsci_d_205_202;
  reg [2:0] chn_data_out_rsci_d_201_199;
  reg [5:0] chn_data_out_rsci_d_198_193;
  reg chn_data_out_rsci_d_192;
  reg chn_data_out_rsci_d_191;
  reg chn_data_out_rsci_d_190;
  reg [3:0] chn_data_out_rsci_d_189_186;
  reg [2:0] chn_data_out_rsci_d_185_183;
  reg [5:0] chn_data_out_rsci_d_182_177;
  reg chn_data_out_rsci_d_176;
  reg chn_data_out_rsci_d_175;
  reg chn_data_out_rsci_d_174;
  reg [3:0] chn_data_out_rsci_d_173_170;
  reg [2:0] chn_data_out_rsci_d_169_167;
  reg [5:0] chn_data_out_rsci_d_166_161;
  reg chn_data_out_rsci_d_160;
  reg chn_data_out_rsci_d_159;
  reg chn_data_out_rsci_d_158;
  reg [3:0] chn_data_out_rsci_d_157_154;
  reg [2:0] chn_data_out_rsci_d_153_151;
  reg [5:0] chn_data_out_rsci_d_150_145;
  reg chn_data_out_rsci_d_144;
  reg chn_data_out_rsci_d_143;
  reg chn_data_out_rsci_d_142;
  reg [3:0] chn_data_out_rsci_d_141_138;
  reg [2:0] chn_data_out_rsci_d_137_135;
  reg [5:0] chn_data_out_rsci_d_134_129;
  reg chn_data_out_rsci_d_128;
  reg chn_data_out_rsci_d_127;
  reg chn_data_out_rsci_d_126;
  reg [3:0] chn_data_out_rsci_d_125_122;
  reg [2:0] chn_data_out_rsci_d_121_119;
  reg [5:0] chn_data_out_rsci_d_118_113;
  reg chn_data_out_rsci_d_112;
  reg chn_data_out_rsci_d_111;
  reg chn_data_out_rsci_d_110;
  reg [3:0] chn_data_out_rsci_d_109_106;
  reg [2:0] chn_data_out_rsci_d_105_103;
  reg [5:0] chn_data_out_rsci_d_102_97;
  reg chn_data_out_rsci_d_96;
  reg chn_data_out_rsci_d_95;
  reg chn_data_out_rsci_d_94;
  reg [3:0] chn_data_out_rsci_d_93_90;
  reg [2:0] chn_data_out_rsci_d_89_87;
  reg [5:0] chn_data_out_rsci_d_86_81;
  reg chn_data_out_rsci_d_80;
  reg chn_data_out_rsci_d_79;
  reg chn_data_out_rsci_d_78;
  reg [3:0] chn_data_out_rsci_d_77_74;
  reg [2:0] chn_data_out_rsci_d_73_71;
  reg [5:0] chn_data_out_rsci_d_70_65;
  reg chn_data_out_rsci_d_64;
  reg chn_data_out_rsci_d_63;
  reg chn_data_out_rsci_d_62;
  reg [3:0] chn_data_out_rsci_d_61_58;
  reg [2:0] chn_data_out_rsci_d_57_55;
  reg [5:0] chn_data_out_rsci_d_54_49;
  reg chn_data_out_rsci_d_48;
  reg chn_data_out_rsci_d_47;
  reg chn_data_out_rsci_d_46;
  reg [3:0] chn_data_out_rsci_d_45_42;
  reg [2:0] chn_data_out_rsci_d_41_39;
  reg [5:0] chn_data_out_rsci_d_38_33;
  reg chn_data_out_rsci_d_32;
  reg chn_data_out_rsci_d_31;
  reg chn_data_out_rsci_d_30;
  reg [3:0] chn_data_out_rsci_d_29_26;
  reg [2:0] chn_data_out_rsci_d_25_23;
  reg [5:0] chn_data_out_rsci_d_22_17;
  reg chn_data_out_rsci_d_16;
  reg chn_data_out_rsci_d_15;
  reg chn_data_out_rsci_d_14;
  reg [3:0] chn_data_out_rsci_d_13_10;
  reg [2:0] chn_data_out_rsci_d_9_7;
  reg [5:0] chn_data_out_rsci_d_6_1;
  reg chn_data_out_rsci_d_0;
  wire [1:0] fsm_output;
  wire IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  wire FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp;
  wire IsDenorm_5U_10U_7_or_3_tmp;
  wire IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  wire FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp;
  wire IsDenorm_5U_10U_7_or_2_tmp;
  wire IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  wire FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp;
  wire IsDenorm_5U_10U_7_or_1_tmp;
  wire IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  wire FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp;
  wire IsDenorm_5U_10U_7_or_tmp;
  wire IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  wire FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp;
  wire IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  wire FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp;
  wire IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
  wire FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp;
  wire IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
  wire FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp;
  wire IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  wire FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp;
  wire IsDenorm_5U_10U_2_or_3_tmp;
  wire IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  wire FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp;
  wire IsDenorm_5U_10U_2_or_2_tmp;
  wire IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  wire FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp;
  wire IsDenorm_5U_10U_2_or_1_tmp;
  wire IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  wire FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp;
  wire IsDenorm_5U_10U_2_or_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  wire FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp;
  wire IsDenorm_5U_10U_1_or_3_tmp;
  wire IsDenorm_5U_10U_or_3_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
  wire FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp;
  wire IsDenorm_5U_10U_1_or_2_tmp;
  wire IsDenorm_5U_10U_or_2_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
  wire FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp;
  wire IsDenorm_5U_10U_1_or_1_tmp;
  wire IsDenorm_5U_10U_or_1_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  wire FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp;
  wire IsDenorm_5U_10U_1_or_tmp;
  wire IsDenorm_5U_10U_or_tmp;
  wire IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp;
  wire IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp;
  wire IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp;
  wire IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp;
  wire m_row3_4_FpMantRNE_23U_11U_3_else_and_tmp;
  wire m_row3_3_FpMantRNE_23U_11U_3_else_and_tmp;
  wire m_row3_2_FpMantRNE_23U_11U_3_else_and_tmp;
  wire m_row3_1_FpMantRNE_23U_11U_3_else_and_tmp;
  wire m_row2_4_FpMantRNE_23U_11U_2_else_and_tmp;
  wire m_row2_3_FpMantRNE_23U_11U_2_else_and_tmp;
  wire m_row2_2_FpMantRNE_23U_11U_2_else_and_tmp;
  wire m_row2_1_FpMantRNE_23U_11U_2_else_and_tmp;
  wire m_row1_4_FpMantRNE_23U_11U_1_else_and_tmp;
  wire m_row1_3_FpMantRNE_23U_11U_1_else_and_tmp;
  wire m_row1_2_FpMantRNE_23U_11U_1_else_and_tmp;
  wire m_row1_1_FpMantRNE_23U_11U_1_else_and_tmp;
  wire m_row0_4_FpMantRNE_23U_11U_else_and_tmp;
  wire m_row0_3_FpMantRNE_23U_11U_else_and_tmp;
  wire m_row0_2_FpMantRNE_23U_11U_else_and_tmp;
  wire m_row0_1_FpMantRNE_23U_11U_else_and_tmp;
  wire o_col3_4_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp;
  wire o_col3_3_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp;
  wire o_col3_2_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp;
  wire o_col3_1_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp;
  wire o_col2_4_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp;
  wire o_col2_3_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp;
  wire o_col2_2_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp;
  wire o_col2_1_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp;
  wire o_col1_4_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp;
  wire o_col1_3_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp;
  wire o_col1_2_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp;
  wire o_col1_1_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp;
  wire o_col0_4_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp;
  wire o_col0_3_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp;
  wire o_col0_2_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp;
  wire o_col0_1_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp;
  wire o_col3_4_FpMantRNE_23U_11U_7_else_and_tmp;
  wire o_col3_3_FpMantRNE_23U_11U_7_else_and_tmp;
  wire o_col3_2_FpMantRNE_23U_11U_7_else_and_tmp;
  wire o_col3_1_FpMantRNE_23U_11U_7_else_and_tmp;
  wire o_col2_4_FpMantRNE_23U_11U_6_else_and_tmp;
  wire o_col2_3_FpMantRNE_23U_11U_6_else_and_tmp;
  wire o_col2_2_FpMantRNE_23U_11U_6_else_and_tmp;
  wire o_col2_1_FpMantRNE_23U_11U_6_else_and_tmp;
  wire o_col1_4_FpMantRNE_23U_11U_5_else_and_tmp;
  wire o_col1_3_FpMantRNE_23U_11U_5_else_and_tmp;
  wire o_col1_2_FpMantRNE_23U_11U_5_else_and_tmp;
  wire o_col1_1_FpMantRNE_23U_11U_5_else_and_tmp;
  wire o_col0_4_FpMantRNE_23U_11U_4_else_and_tmp;
  wire o_col0_3_FpMantRNE_23U_11U_4_else_and_tmp;
  wire o_col0_2_FpMantRNE_23U_11U_4_else_and_tmp;
  wire o_col0_1_FpMantRNE_23U_11U_4_else_and_tmp;
  wire IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp;
  wire IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp;
  wire IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_tmp;
  wire IsNaN_6U_10U_16_nor_15_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_14_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_13_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_tmp;
  wire IsNaN_6U_10U_16_nor_12_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_11_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_10_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_9_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_8_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_7_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_6_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_5_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_4_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_3_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_2_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_1_tmp;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_tmp;
  wire IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp;
  wire IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_3_tmp;
  wire IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_2_tmp;
  wire IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_1_tmp;
  wire IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_tmp;
  wire IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp;
  wire IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp;
  wire IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp;
  wire IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp;
  wire IsNaN_6U_10U_10_nor_1_tmp;
  wire IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp;
  wire IsNaN_6U_10U_9_nor_3_tmp;
  wire IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp;
  wire IsNaN_6U_10U_9_nor_2_tmp;
  wire IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp;
  wire IsNaN_6U_10U_9_nor_1_tmp;
  wire IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp;
  wire and_dcpl_3;
  wire and_dcpl_52;
  wire or_dcpl_1;
  wire and_dcpl_57;
  wire not_tmp_35;
  wire or_tmp_5;
  wire or_tmp_8;
  wire nand_tmp_2;
  wire or_tmp_16;
  wire or_tmp_19;
  wire or_tmp_22;
  wire or_tmp_25;
  wire nand_tmp_15;
  wire or_tmp_27;
  wire nand_tmp_16;
  wire or_tmp_30;
  wire or_tmp_33;
  wire or_tmp_36;
  wire or_tmp_39;
  wire or_tmp_42;
  wire nand_tmp_31;
  wire or_tmp_44;
  wire or_tmp_45;
  wire and_tmp_1;
  wire mux_tmp_35;
  wire or_tmp_48;
  wire or_tmp_52;
  wire or_tmp_57;
  wire or_tmp_65;
  wire mux_tmp_49;
  wire mux_tmp_51;
  wire not_tmp_81;
  wire mux_tmp_56;
  wire not_tmp_83;
  wire mux_tmp_61;
  wire not_tmp_85;
  wire mux_tmp_69;
  wire not_tmp_90;
  wire nor_tmp_72;
  wire mux_tmp_73;
  wire not_tmp_92;
  wire mux_tmp_76;
  wire mux_tmp_81;
  wire not_tmp_96;
  wire nor_tmp_78;
  wire mux_tmp_85;
  wire not_tmp_98;
  wire mux_tmp_88;
  wire mux_tmp_93;
  wire not_tmp_102;
  wire nor_tmp_84;
  wire mux_tmp_97;
  wire not_tmp_104;
  wire mux_tmp_100;
  wire or_tmp_170;
  wire not_tmp_109;
  wire or_tmp_183;
  wire not_tmp_112;
  wire or_tmp_196;
  wire not_tmp_115;
  wire or_tmp_211;
  wire not_tmp_120;
  wire mux_tmp_142;
  wire or_tmp_224;
  wire not_tmp_123;
  wire mux_tmp_151;
  wire nor_tmp_118;
  wire or_tmp_243;
  wire not_tmp_128;
  wire mux_tmp_162;
  wire nor_tmp_127;
  wire mux_tmp_169;
  wire not_tmp_134;
  wire mux_tmp_172;
  wire nor_tmp_130;
  wire mux_tmp_176;
  wire not_tmp_138;
  wire mux_tmp_179;
  wire nor_tmp_133;
  wire mux_tmp_183;
  wire not_tmp_142;
  wire mux_tmp_186;
  wire mux_tmp_191;
  wire mux_tmp_192;
  wire mux_tmp_193;
  wire not_tmp_148;
  wire or_tmp_286;
  wire mux_tmp_198;
  wire or_tmp_287;
  wire or_tmp_288;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire or_tmp_290;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire mux_tmp_204;
  wire mux_tmp_205;
  wire mux_tmp_206;
  wire mux_tmp_207;
  wire mux_tmp_208;
  wire mux_tmp_212;
  wire or_tmp_302;
  wire or_tmp_303;
  wire mux_tmp_219;
  wire or_tmp_319;
  wire or_tmp_320;
  wire mux_tmp_228;
  wire or_tmp_336;
  wire or_tmp_337;
  wire mux_tmp_237;
  wire mux_tmp_246;
  wire mux_tmp_250;
  wire mux_tmp_254;
  wire or_tmp_359;
  wire or_tmp_360;
  wire mux_tmp_258;
  wire or_tmp_376;
  wire or_tmp_377;
  wire mux_tmp_267;
  wire or_tmp_393;
  wire or_tmp_394;
  wire mux_tmp_276;
  wire mux_tmp_291;
  wire or_tmp_419;
  wire or_tmp_420;
  wire mux_tmp_299;
  wire or_tmp_437;
  wire mux_tmp_308;
  wire mux_tmp_311;
  wire mux_tmp_313;
  wire or_tmp_438;
  wire or_tmp_441;
  wire or_tmp_442;
  wire mux_tmp_317;
  wire mux_tmp_329;
  wire or_tmp_465;
  wire or_tmp_466;
  wire mux_tmp_340;
  wire mux_tmp_351;
  wire or_tmp_485;
  wire or_tmp_486;
  wire mux_tmp_355;
  wire mux_tmp_364;
  wire or_tmp_510;
  wire or_tmp_513;
  wire or_tmp_514;
  wire mux_tmp_371;
  wire mux_tmp_380;
  wire or_tmp_532;
  wire or_tmp_533;
  wire mux_tmp_384;
  wire mux_tmp_393;
  wire or_tmp_551;
  wire or_tmp_552;
  wire mux_tmp_397;
  wire or_tmp_576;
  wire or_tmp_579;
  wire or_tmp_580;
  wire mux_tmp_413;
  wire nand_tmp_61;
  wire mux_tmp_429;
  wire not_tmp_203;
  wire mux_tmp_435;
  wire not_tmp_204;
  wire or_tmp_614;
  wire not_tmp_205;
  wire mux_tmp_443;
  wire or_tmp_624;
  wire not_tmp_208;
  wire or_tmp_634;
  wire not_tmp_211;
  wire mux_tmp_457;
  wire or_tmp_640;
  wire not_tmp_212;
  wire mux_tmp_460;
  wire and_tmp_56;
  wire or_tmp_721;
  wire or_tmp_723;
  wire or_tmp_736;
  wire or_tmp_738;
  wire or_tmp_751;
  wire or_tmp_753;
  wire or_tmp_774;
  wire or_tmp_823;
  wire mux_tmp_570;
  wire or_tmp_828;
  wire mux_tmp_603;
  wire or_tmp_923;
  wire mux_tmp_622;
  wire or_tmp_963;
  wire or_tmp_966;
  wire or_tmp_976;
  wire or_tmp_977;
  wire and_dcpl_64;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire or_dcpl_21;
  wire or_dcpl_23;
  wire and_dcpl_74;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_81;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire or_dcpl_64;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_99;
  wire and_dcpl_101;
  wire or_dcpl_69;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire or_dcpl_70;
  wire and_dcpl_110;
  wire and_dcpl_112;
  wire and_dcpl_117;
  wire or_dcpl_75;
  wire and_dcpl_120;
  wire and_dcpl_122;
  wire and_dcpl_124;
  wire and_dcpl_129;
  wire or_dcpl_80;
  wire and_dcpl_132;
  wire and_dcpl_134;
  wire and_dcpl_140;
  wire and_dcpl_142;
  wire and_dcpl_147;
  wire or_dcpl_86;
  wire and_dcpl_150;
  wire and_dcpl_152;
  wire and_dcpl_154;
  wire and_dcpl_159;
  wire and_dcpl_161;
  wire or_dcpl_91;
  wire and_dcpl_162;
  wire and_dcpl_164;
  wire or_dcpl_92;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire or_dcpl_93;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire or_dcpl_94;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire or_dcpl_95;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_213;
  wire and_dcpl_214;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire or_dcpl_99;
  wire and_dcpl_231;
  wire and_dcpl_232;
  wire or_dcpl_100;
  wire and_dcpl_238;
  wire and_dcpl_239;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_248;
  wire and_dcpl_253;
  wire or_dcpl_106;
  wire and_dcpl_256;
  wire and_dcpl_259;
  wire and_dcpl_264;
  wire or_dcpl_111;
  wire and_dcpl_267;
  wire and_dcpl_269;
  wire and_dcpl_270;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_279;
  wire and_dcpl_281;
  wire or_dcpl_116;
  wire and_dcpl_282;
  wire and_dcpl_285;
  wire and_dcpl_290;
  wire or_dcpl_121;
  wire and_dcpl_293;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_297;
  wire and_dcpl_298;
  wire and_dcpl_300;
  wire and_dcpl_305;
  wire and_dcpl_307;
  wire or_dcpl_126;
  wire and_dcpl_308;
  wire and_dcpl_311;
  wire and_dcpl_316;
  wire or_dcpl_131;
  wire and_dcpl_319;
  wire and_dcpl_321;
  wire and_dcpl_322;
  wire and_dcpl_323;
  wire and_dcpl_324;
  wire and_dcpl_333;
  wire and_dcpl_334;
  wire and_dcpl_343;
  wire and_dcpl_344;
  wire and_dcpl_353;
  wire and_dcpl_354;
  wire and_dcpl_357;
  wire and_dcpl_363;
  wire and_dcpl_364;
  wire and_dcpl_366;
  wire and_dcpl_369;
  wire and_dcpl_375;
  wire and_dcpl_376;
  wire and_dcpl_378;
  wire and_dcpl_381;
  wire and_dcpl_387;
  wire and_dcpl_388;
  wire mux_tmp_656;
  wire and_dcpl_391;
  wire mux_tmp_657;
  wire and_dcpl_394;
  wire mux_tmp_658;
  wire and_dcpl_397;
  wire or_dcpl_168;
  wire and_dcpl_449;
  wire or_dcpl_170;
  wire and_dcpl_453;
  wire or_dcpl_172;
  wire and_dcpl_457;
  wire or_dcpl_174;
  wire and_dcpl_461;
  wire or_dcpl_176;
  wire and_dcpl_465;
  wire or_dcpl_178;
  wire and_dcpl_469;
  wire or_dcpl_180;
  wire and_dcpl_473;
  wire or_dcpl_182;
  wire and_dcpl_477;
  wire or_dcpl_184;
  wire and_dcpl_481;
  wire or_dcpl_186;
  wire and_dcpl_485;
  wire or_dcpl_188;
  wire and_dcpl_489;
  wire or_dcpl_190;
  wire and_dcpl_493;
  wire or_dcpl_192;
  wire and_dcpl_497;
  wire or_dcpl_194;
  wire and_dcpl_501;
  wire or_dcpl_196;
  wire and_dcpl_505;
  wire or_dcpl_198;
  wire and_dcpl_509;
  wire or_dcpl_200;
  wire or_dcpl_203;
  wire or_dcpl_206;
  wire or_dcpl_209;
  wire or_dcpl_212;
  wire or_dcpl_215;
  wire or_dcpl_218;
  wire or_dcpl_221;
  wire or_dcpl_224;
  wire or_dcpl_227;
  wire or_dcpl_230;
  wire or_dcpl_233;
  wire or_dcpl_236;
  wire or_dcpl_239;
  wire or_dcpl_242;
  wire or_dcpl_245;
  wire or_dcpl_248;
  wire or_dcpl_251;
  wire or_dcpl_254;
  wire or_dcpl_257;
  wire or_dcpl_260;
  wire or_dcpl_263;
  wire or_dcpl_266;
  wire or_dcpl_269;
  wire or_dcpl_272;
  wire or_dcpl_275;
  wire or_dcpl_278;
  wire or_dcpl_281;
  wire or_dcpl_284;
  wire or_dcpl_287;
  wire or_dcpl_290;
  wire or_dcpl_293;
  wire and_dcpl_547;
  wire or_dcpl_296;
  wire or_dcpl_301;
  wire or_dcpl_302;
  wire and_dcpl_644;
  wire and_dcpl_645;
  wire and_dcpl_651;
  wire or_dcpl_303;
  wire and_dcpl_658;
  wire and_dcpl_659;
  wire and_dcpl_665;
  wire and_dcpl_672;
  wire and_dcpl_673;
  wire and_dcpl_679;
  wire and_dcpl_686;
  wire and_dcpl_687;
  wire and_dcpl_693;
  wire and_dcpl_701;
  wire and_dcpl_707;
  wire and_dcpl_715;
  wire and_dcpl_721;
  wire and_dcpl_729;
  wire and_dcpl_735;
  wire and_dcpl_742;
  wire and_dcpl_743;
  wire and_dcpl_749;
  wire and_dcpl_756;
  wire and_dcpl_757;
  wire and_dcpl_763;
  wire and_dcpl_770;
  wire and_dcpl_771;
  wire and_dcpl_777;
  wire and_dcpl_785;
  wire and_dcpl_791;
  wire and_dcpl_799;
  wire and_dcpl_805;
  wire and_dcpl_817;
  wire and_dcpl_823;
  wire and_dcpl_824;
  wire and_dcpl_833;
  wire and_dcpl_834;
  wire and_dcpl_843;
  wire and_dcpl_844;
  wire and_dcpl_853;
  wire and_dcpl_854;
  wire and_dcpl_863;
  wire and_dcpl_864;
  wire and_dcpl_873;
  wire and_dcpl_874;
  wire and_dcpl_883;
  wire and_dcpl_884;
  wire and_dcpl_893;
  wire and_dcpl_894;
  wire and_dcpl_903;
  wire and_dcpl_904;
  wire and_dcpl_913;
  wire and_dcpl_914;
  wire and_dcpl_923;
  wire and_dcpl_924;
  wire and_dcpl_933;
  wire and_dcpl_934;
  wire and_dcpl_943;
  wire and_dcpl_944;
  wire and_dcpl_953;
  wire and_dcpl_954;
  wire and_dcpl_963;
  wire and_dcpl_964;
  wire and_dcpl_973;
  wire and_dcpl_974;
  wire and_dcpl_975;
  wire and_dcpl_977;
  wire and_dcpl_982;
  wire or_dcpl_336;
  wire and_dcpl_985;
  wire and_dcpl_987;
  wire and_dcpl_989;
  wire and_dcpl_994;
  wire and_dcpl_996;
  wire or_dcpl_341;
  wire and_dcpl_997;
  wire and_dcpl_999;
  wire or_dcpl_342;
  wire and_dcpl_1001;
  wire and_dcpl_1002;
  wire or_dcpl_343;
  wire and_dcpl_1004;
  wire and_dcpl_1005;
  wire and_dcpl_1007;
  wire and_dcpl_1008;
  wire or_dcpl_345;
  wire and_dcpl_1010;
  wire and_dcpl_1012;
  wire and_dcpl_1017;
  wire and_dcpl_1019;
  wire or_dcpl_350;
  wire and_dcpl_1020;
  wire and_dcpl_1023;
  wire and_dcpl_1028;
  wire or_dcpl_355;
  wire and_dcpl_1031;
  wire and_dcpl_1033;
  wire and_dcpl_1034;
  wire and_dcpl_1035;
  wire and_dcpl_1036;
  wire and_dcpl_1045;
  wire and_dcpl_1046;
  wire and_dcpl_1049;
  wire and_dcpl_1055;
  wire and_dcpl_1056;
  wire mux_tmp_661;
  wire and_dcpl_1059;
  wire and_dcpl_1061;
  wire and_dcpl_1067;
  wire and_dcpl_1074;
  wire and_dcpl_1075;
  wire and_dcpl_1081;
  wire and_dcpl_1089;
  wire and_dcpl_1095;
  wire and_dcpl_1102;
  wire and_dcpl_1103;
  wire and_dcpl_1109;
  wire and_dcpl_1119;
  wire and_dcpl_1122;
  wire or_dcpl_366;
  wire and_dcpl_1126;
  wire or_dcpl_367;
  wire and_dcpl_1129;
  wire and_dcpl_1131;
  wire and_dcpl_1133;
  wire and_dcpl_1136;
  wire and_dcpl_1138;
  wire and_dcpl_1141;
  wire and_dcpl_1143;
  wire and_dcpl_1146;
  wire and_dcpl_1148;
  wire and_dcpl_1151;
  wire and_dcpl_1153;
  wire and_dcpl_1156;
  wire and_dcpl_1158;
  wire and_dcpl_1161;
  wire and_dcpl_1163;
  wire and_dcpl_1166;
  wire and_dcpl_1168;
  wire and_dcpl_1171;
  wire and_dcpl_1173;
  wire and_dcpl_1176;
  wire and_dcpl_1178;
  wire and_dcpl_1181;
  wire and_dcpl_1183;
  wire and_dcpl_1186;
  wire and_dcpl_1188;
  wire and_dcpl_1191;
  wire and_dcpl_1193;
  wire and_dcpl_1196;
  wire and_dcpl_1198;
  wire and_dcpl_1201;
  wire and_dcpl_1203;
  wire and_dcpl_1206;
  wire and_dcpl_1208;
  wire or_dcpl_368;
  wire or_tmp_1099;
  reg [5:0] FpAdd_6U_10U_4_o_expo_1_lpi_2;
  reg [9:0] FpAdd_6U_10U_4_o_mant_1_lpi_2;
  reg [5:0] FpAdd_6U_10U_4_o_expo_2_lpi_2;
  reg [9:0] FpAdd_6U_10U_4_o_mant_2_lpi_2;
  reg [5:0] FpAdd_6U_10U_4_o_expo_3_lpi_2;
  reg [9:0] FpAdd_6U_10U_4_o_mant_3_lpi_2;
  reg [5:0] FpAdd_6U_10U_4_o_expo_lpi_2;
  reg [9:0] FpAdd_6U_10U_4_o_mant_lpi_2;
  reg [5:0] FpAdd_6U_10U_5_o_expo_1_lpi_2;
  reg [9:0] FpAdd_6U_10U_5_o_mant_1_lpi_2;
  reg [5:0] FpAdd_6U_10U_5_o_expo_2_lpi_2;
  reg [9:0] FpAdd_6U_10U_5_o_mant_2_lpi_2;
  reg [5:0] FpAdd_6U_10U_5_o_expo_3_lpi_2;
  reg [9:0] FpAdd_6U_10U_5_o_mant_3_lpi_2;
  reg [5:0] FpAdd_6U_10U_5_o_expo_lpi_2;
  reg [9:0] FpAdd_6U_10U_5_o_mant_lpi_2;
  reg [5:0] FpAdd_6U_10U_6_o_expo_1_lpi_2;
  reg [9:0] FpAdd_6U_10U_6_o_mant_1_lpi_2;
  reg [5:0] FpAdd_6U_10U_6_o_expo_2_lpi_2;
  reg [9:0] FpAdd_6U_10U_6_o_mant_2_lpi_2;
  reg [5:0] FpAdd_6U_10U_6_o_expo_3_lpi_2;
  reg [9:0] FpAdd_6U_10U_6_o_mant_3_lpi_2;
  reg [5:0] FpAdd_6U_10U_6_o_expo_lpi_2;
  reg [9:0] FpAdd_6U_10U_6_o_mant_lpi_2;
  reg [5:0] FpAdd_6U_10U_7_o_expo_1_lpi_2;
  reg [9:0] FpAdd_6U_10U_7_o_mant_1_lpi_2;
  reg [5:0] FpAdd_6U_10U_7_o_expo_2_lpi_2;
  reg [9:0] FpAdd_6U_10U_7_o_mant_2_lpi_2;
  reg [5:0] FpAdd_6U_10U_7_o_expo_3_lpi_2;
  reg [9:0] FpAdd_6U_10U_7_o_mant_3_lpi_2;
  reg [5:0] FpAdd_6U_10U_7_o_expo_lpi_2;
  reg [9:0] FpAdd_6U_10U_7_o_mant_lpi_2;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_6;
  reg FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_1_sva;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_1_sva;
  reg IsNaN_6U_10U_land_1_lpi_1_dfm;
  reg IsNaN_6U_10U_1_land_1_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_6;
  reg FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_2_sva;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_2_sva;
  reg IsNaN_6U_10U_land_2_lpi_1_dfm;
  reg IsNaN_6U_10U_1_land_2_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_6;
  reg FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_3_sva;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_3_sva;
  reg IsNaN_6U_10U_land_3_lpi_1_dfm;
  reg IsNaN_6U_10U_1_land_3_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_6;
  reg FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_qr_3_0_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_sva;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_sva;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm;
  reg [9:0] FpAdd_6U_10U_o_mant_lpi_1_dfm_2;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_6;
  reg FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_1_sva;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_1_sva;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm;
  reg IsNaN_6U_10U_3_land_1_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_6;
  reg FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_2_sva;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_2_sva;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm;
  reg IsNaN_6U_10U_3_land_2_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_6;
  reg FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_3_sva;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_3_sva;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm;
  reg IsNaN_6U_10U_3_land_3_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_6;
  reg FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_sva;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_sva;
  reg IsNaN_6U_10U_3_land_lpi_1_dfm;
  reg [9:0] FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_6;
  reg FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_1_sva;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_1_sva;
  reg IsNaN_6U_10U_4_land_1_lpi_1_dfm;
  reg IsNaN_6U_10U_5_land_1_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_6;
  reg FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_2_sva;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_2_sva;
  reg IsNaN_6U_10U_4_land_2_lpi_1_dfm;
  reg IsNaN_6U_10U_5_land_2_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_6;
  reg FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_3_sva;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_3_sva;
  reg IsNaN_6U_10U_4_land_3_lpi_1_dfm;
  reg IsNaN_6U_10U_5_land_3_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_6;
  reg FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_sva;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_sva;
  reg IsNaN_6U_10U_5_land_lpi_1_dfm;
  reg [9:0] FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_1_sva;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_1_sva;
  reg IsNaN_6U_10U_6_land_1_lpi_1_dfm;
  reg IsNaN_6U_10U_7_land_1_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_2_sva;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_2_sva;
  reg IsNaN_6U_10U_6_land_2_lpi_1_dfm;
  reg IsNaN_6U_10U_7_land_2_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_3_sva;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_3_sva;
  reg IsNaN_6U_10U_6_land_3_lpi_1_dfm;
  reg IsNaN_6U_10U_7_land_3_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_6;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_6;
  reg [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_1;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_sva;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_sva;
  reg IsNaN_6U_10U_7_land_lpi_1_dfm;
  reg [9:0] FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2;
  reg [16:0] m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva;
  reg [16:0] m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva;
  reg [16:0] m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva;
  reg [16:0] m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva;
  reg [16:0] m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva;
  reg [16:0] m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva;
  reg [16:0] m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva;
  reg [16:0] m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva;
  reg FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2;
  reg FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2;
  reg FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2;
  reg FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2;
  reg data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs;
  reg data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg IsNaN_6U_10U_16_land_1_lpi_1_dfm_3;
  reg data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_2_lpi_1_dfm_3;
  reg data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_3_lpi_1_dfm_3;
  reg data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_4_lpi_1_dfm_3;
  reg data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_5_lpi_1_dfm_3;
  reg data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_6_lpi_1_dfm_3;
  reg data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_7_lpi_1_dfm_3;
  reg data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_8_lpi_1_dfm_3;
  reg data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_9_lpi_1_dfm_3;
  reg data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_10_lpi_1_dfm_3;
  reg data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_11_lpi_1_dfm_3;
  reg data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_12_lpi_1_dfm_3;
  reg data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_14_lpi_1_dfm_3;
  reg data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg IsNaN_6U_10U_16_land_15_lpi_1_dfm_3;
  reg data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  reg FpAdd_6U_10U_2_o_sign_lpi_1_dfm_4;
  reg FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_o_sign_lpi_1_dfm_4;
  reg FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5;
  reg FpAdd_6U_10U_o_sign_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5;
  reg IsNaN_6U_10U_14_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_14_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_14_land_1_lpi_1_dfm_5;
  reg [9:0] FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7;
  reg IsNaN_6U_10U_12_land_3_lpi_1_dfm_4;
  reg FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_4;
  reg FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_12_land_2_lpi_1_dfm_4;
  reg FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_4;
  reg FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_12_land_1_lpi_1_dfm_4;
  reg FpAdd_6U_10U_o_sign_3_lpi_1_dfm_4;
  reg [9:0] FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7;
  reg IsNaN_6U_10U_10_land_3_lpi_1_dfm_4;
  reg IsNaN_6U_10U_10_land_3_lpi_1_dfm_5;
  reg FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_4;
  reg FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_10_land_2_lpi_1_dfm_4;
  reg IsNaN_6U_10U_10_land_2_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_4;
  reg FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_10_land_1_lpi_1_dfm_4;
  reg IsNaN_6U_10U_10_land_1_lpi_1_dfm_5;
  reg FpAdd_6U_10U_o_sign_2_lpi_1_dfm_4;
  reg [9:0] FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_7;
  reg [9:0] FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_o_mant_1_lpi_1_dfm_7;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_5;
  reg FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_4;
  reg FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_4;
  reg FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_8_land_1_lpi_1_dfm_4;
  reg IsNaN_6U_10U_8_land_1_lpi_1_dfm_5;
  reg FpAdd_6U_10U_o_sign_1_lpi_1_dfm_4;
  reg IsNaN_6U_10U_14_land_lpi_1_dfm_5;
  reg [9:0] FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7;
  reg IsNaN_6U_10U_12_land_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5;
  reg [9:0] FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7;
  reg IsNaN_6U_10U_10_land_lpi_1_dfm_4;
  reg IsNaN_6U_10U_10_land_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5;
  reg [9:0] FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_7;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_5;
  reg FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_4;
  reg FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_15_land_lpi_1_dfm_4;
  reg IsNaN_6U_10U_15_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_15_land_3_lpi_1_dfm_4;
  reg IsNaN_6U_10U_15_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_15_land_2_lpi_1_dfm_4;
  reg IsNaN_6U_10U_15_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_15_land_1_lpi_1_dfm_4;
  reg IsNaN_6U_10U_15_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_13_land_lpi_1_dfm_4;
  reg IsNaN_6U_10U_13_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_13_land_3_lpi_1_dfm_4;
  reg IsNaN_6U_10U_13_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_13_land_2_lpi_1_dfm_3;
  reg IsNaN_6U_10U_13_land_1_lpi_1_dfm_4;
  reg IsNaN_6U_10U_13_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_11_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_11_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_11_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_9_land_lpi_1_dfm_3;
  reg IsNaN_6U_10U_9_land_3_lpi_1_dfm_3;
  reg IsNaN_6U_10U_9_land_2_lpi_1_dfm_3;
  reg IsNaN_6U_10U_9_land_1_lpi_1_dfm_5;
  reg [5:0] o_data_data_15_6_1_sva_7;
  reg [5:0] o_data_data_15_6_1_sva_8;
  reg [5:0] o_data_data_14_6_1_sva_7;
  reg [5:0] o_data_data_14_6_1_sva_8;
  reg [5:0] o_data_data_13_6_1_sva_7;
  reg [5:0] o_data_data_13_6_1_sva_8;
  reg [5:0] o_data_data_12_6_1_sva_7;
  reg [5:0] o_data_data_12_6_1_sva_8;
  reg [5:0] o_data_data_11_6_1_sva_7;
  reg [5:0] o_data_data_11_6_1_sva_8;
  reg [5:0] o_data_data_10_6_1_sva_7;
  reg [5:0] o_data_data_10_6_1_sva_8;
  reg [5:0] o_data_data_9_6_1_sva_7;
  reg [5:0] o_data_data_9_6_1_sva_8;
  reg [5:0] o_data_data_8_6_1_sva_7;
  reg [5:0] o_data_data_8_6_1_sva_8;
  reg [5:0] o_data_data_7_6_1_sva_7;
  reg [5:0] o_data_data_7_6_1_sva_8;
  reg [5:0] o_data_data_6_6_1_sva_7;
  reg [5:0] o_data_data_6_6_1_sva_8;
  reg [5:0] o_data_data_5_6_1_sva_7;
  reg [5:0] o_data_data_5_6_1_sva_8;
  reg [5:0] o_data_data_4_6_1_sva_7;
  reg [5:0] o_data_data_4_6_1_sva_8;
  reg [5:0] o_data_data_3_6_1_sva_7;
  reg [5:0] o_data_data_3_6_1_sva_8;
  reg [5:0] o_data_data_2_6_1_sva_7;
  reg [5:0] o_data_data_2_6_1_sva_8;
  reg [5:0] o_data_data_1_6_1_sva_7;
  reg [5:0] o_data_data_1_6_1_sva_8;
  reg [5:0] o_data_data_0_6_1_sva_7;
  reg [5:0] o_data_data_0_6_1_sva_8;
  reg [5:0] o_data_data_15_6_1_sva_9;
  reg [5:0] o_data_data_15_6_1_sva_10;
  reg [3:0] o_data_data_15_13_10_sva_5;
  reg [3:0] o_data_data_15_13_10_sva_6;
  reg [2:0] o_data_data_15_9_7_sva_5;
  reg [2:0] o_data_data_15_9_7_sva_6;
  reg [5:0] o_data_data_14_6_1_sva_9;
  reg [5:0] o_data_data_14_6_1_sva_10;
  reg [3:0] o_data_data_14_13_10_sva_5;
  reg [3:0] o_data_data_14_13_10_sva_6;
  reg [2:0] o_data_data_14_9_7_sva_5;
  reg [2:0] o_data_data_14_9_7_sva_6;
  reg [5:0] o_data_data_13_6_1_sva_9;
  reg [5:0] o_data_data_13_6_1_sva_10;
  reg [3:0] o_data_data_13_13_10_sva_5;
  reg [3:0] o_data_data_13_13_10_sva_6;
  reg [2:0] o_data_data_13_9_7_sva_5;
  reg [2:0] o_data_data_13_9_7_sva_6;
  reg [5:0] o_data_data_12_6_1_sva_9;
  reg [5:0] o_data_data_12_6_1_sva_10;
  reg [3:0] o_data_data_12_13_10_sva_5;
  reg [3:0] o_data_data_12_13_10_sva_6;
  reg [2:0] o_data_data_12_9_7_sva_5;
  reg [2:0] o_data_data_12_9_7_sva_6;
  reg [5:0] o_data_data_11_6_1_sva_9;
  reg [5:0] o_data_data_11_6_1_sva_10;
  reg [3:0] o_data_data_11_13_10_sva_5;
  reg [3:0] o_data_data_11_13_10_sva_6;
  reg [2:0] o_data_data_11_9_7_sva_5;
  reg [2:0] o_data_data_11_9_7_sva_6;
  reg [5:0] o_data_data_10_6_1_sva_9;
  reg [5:0] o_data_data_10_6_1_sva_10;
  reg [3:0] o_data_data_10_13_10_sva_5;
  reg [3:0] o_data_data_10_13_10_sva_6;
  reg [2:0] o_data_data_10_9_7_sva_5;
  reg [2:0] o_data_data_10_9_7_sva_6;
  reg [5:0] o_data_data_9_6_1_sva_9;
  reg [5:0] o_data_data_9_6_1_sva_10;
  reg [3:0] o_data_data_9_13_10_sva_5;
  reg [3:0] o_data_data_9_13_10_sva_6;
  reg [2:0] o_data_data_9_9_7_sva_5;
  reg [2:0] o_data_data_9_9_7_sva_6;
  reg [5:0] o_data_data_8_6_1_sva_9;
  reg [5:0] o_data_data_8_6_1_sva_10;
  reg [3:0] o_data_data_8_13_10_sva_5;
  reg [3:0] o_data_data_8_13_10_sva_6;
  reg [2:0] o_data_data_8_9_7_sva_5;
  reg [2:0] o_data_data_8_9_7_sva_6;
  reg [5:0] o_data_data_7_6_1_sva_9;
  reg [5:0] o_data_data_7_6_1_sva_10;
  reg [3:0] o_data_data_7_13_10_sva_5;
  reg [3:0] o_data_data_7_13_10_sva_6;
  reg [2:0] o_data_data_7_9_7_sva_5;
  reg [2:0] o_data_data_7_9_7_sva_6;
  reg [5:0] o_data_data_6_6_1_sva_9;
  reg [5:0] o_data_data_6_6_1_sva_10;
  reg [3:0] o_data_data_6_13_10_sva_5;
  reg [3:0] o_data_data_6_13_10_sva_6;
  reg [2:0] o_data_data_6_9_7_sva_5;
  reg [2:0] o_data_data_6_9_7_sva_6;
  reg [5:0] o_data_data_5_6_1_sva_9;
  reg [5:0] o_data_data_5_6_1_sva_10;
  reg [3:0] o_data_data_5_13_10_sva_5;
  reg [3:0] o_data_data_5_13_10_sva_6;
  reg [2:0] o_data_data_5_9_7_sva_5;
  reg [2:0] o_data_data_5_9_7_sva_6;
  reg [5:0] o_data_data_4_6_1_sva_9;
  reg [5:0] o_data_data_4_6_1_sva_10;
  reg [3:0] o_data_data_4_13_10_sva_5;
  reg [3:0] o_data_data_4_13_10_sva_6;
  reg [2:0] o_data_data_4_9_7_sva_5;
  reg [2:0] o_data_data_4_9_7_sva_6;
  reg [5:0] o_data_data_3_6_1_sva_9;
  reg [5:0] o_data_data_3_6_1_sva_10;
  reg [3:0] o_data_data_3_13_10_sva_5;
  reg [3:0] o_data_data_3_13_10_sva_6;
  reg [2:0] o_data_data_3_9_7_sva_5;
  reg [2:0] o_data_data_3_9_7_sva_6;
  reg [5:0] o_data_data_2_6_1_sva_9;
  reg [5:0] o_data_data_2_6_1_sva_10;
  reg [3:0] o_data_data_2_13_10_sva_5;
  reg [3:0] o_data_data_2_13_10_sva_6;
  reg [2:0] o_data_data_2_9_7_sva_5;
  reg [2:0] o_data_data_2_9_7_sva_6;
  reg [5:0] o_data_data_1_6_1_sva_9;
  reg [5:0] o_data_data_1_6_1_sva_10;
  reg [3:0] o_data_data_1_13_10_sva_5;
  reg [3:0] o_data_data_1_13_10_sva_6;
  reg [2:0] o_data_data_1_9_7_sva_5;
  reg [2:0] o_data_data_1_9_7_sva_6;
  reg [5:0] o_data_data_0_6_1_sva_9;
  reg [5:0] o_data_data_0_6_1_sva_10;
  reg [3:0] o_data_data_0_13_10_sva_5;
  reg [3:0] o_data_data_0_13_10_sva_6;
  reg [2:0] o_data_data_0_9_7_sva_5;
  reg [2:0] o_data_data_0_9_7_sva_6;
  reg [23:0] FpAdd_6U_10U_7_int_mant_p1_sva_3;
  reg [23:0] FpAdd_6U_10U_7_int_mant_p1_3_sva_3;
  reg [23:0] FpAdd_6U_10U_7_int_mant_p1_2_sva_3;
  reg [23:0] FpAdd_6U_10U_7_int_mant_p1_1_sva_3;
  reg [23:0] FpAdd_6U_10U_6_int_mant_p1_sva_3;
  reg [23:0] FpAdd_6U_10U_6_int_mant_p1_3_sva_3;
  reg [23:0] FpAdd_6U_10U_6_int_mant_p1_2_sva_3;
  reg [23:0] FpAdd_6U_10U_6_int_mant_p1_1_sva_3;
  reg [23:0] FpAdd_6U_10U_5_int_mant_p1_sva_3;
  reg [23:0] FpAdd_6U_10U_5_int_mant_p1_3_sva_3;
  reg [23:0] FpAdd_6U_10U_5_int_mant_p1_2_sva_3;
  reg [23:0] FpAdd_6U_10U_5_int_mant_p1_1_sva_3;
  reg [23:0] FpAdd_6U_10U_4_int_mant_p1_sva_3;
  reg [23:0] FpAdd_6U_10U_4_int_mant_p1_3_sva_3;
  reg [23:0] FpAdd_6U_10U_4_int_mant_p1_2_sva_3;
  reg [23:0] FpAdd_6U_10U_4_int_mant_p1_1_sva_3;
  reg m_row0_unequal_tmp_3;
  reg m_row0_unequal_tmp_4;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_7;
  reg FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_1_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_1_sva_2;
  reg IsNaN_6U_10U_1_land_1_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_7;
  reg FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_2_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_2_sva_2;
  reg IsNaN_6U_10U_1_land_2_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_7;
  reg FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_3_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_3_sva_2;
  reg IsNaN_6U_10U_1_land_3_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_7;
  reg FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_sva_2;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_3;
  reg [9:0] FpAdd_6U_10U_o_mant_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_o_mant_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_7;
  reg FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_1_sva_2;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_3;
  reg IsNaN_6U_10U_3_land_1_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_7;
  reg FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_2_sva_2;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_3;
  reg IsNaN_6U_10U_3_land_2_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_7;
  reg FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_3_sva_2;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_3;
  reg IsNaN_6U_10U_3_land_3_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_7;
  reg FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_1_a_int_mant_p1_sva_2;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_sva_2;
  reg IsNaN_6U_10U_3_land_lpi_1_dfm_3;
  reg [9:0] FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_1_o_mant_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_7;
  reg FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_1_sva_2;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_1_sva_2;
  reg IsNaN_6U_10U_4_land_1_lpi_1_dfm_3;
  reg IsNaN_6U_10U_5_land_1_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_7;
  reg FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_2_sva_2;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_2_sva_2;
  reg IsNaN_6U_10U_4_land_2_lpi_1_dfm_3;
  reg IsNaN_6U_10U_5_land_2_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_7;
  reg FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_3_sva_2;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_3_sva_2;
  reg IsNaN_6U_10U_4_land_3_lpi_1_dfm_3;
  reg IsNaN_6U_10U_5_land_3_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_7;
  reg FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_2_a_int_mant_p1_sva_2;
  reg [22:0] FpAdd_6U_10U_2_b_int_mant_p1_sva_2;
  reg IsNaN_6U_10U_5_land_lpi_1_dfm_3;
  reg [9:0] FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_2_o_mant_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_7;
  reg FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_1_sva_2;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_1_sva_2;
  reg IsNaN_6U_10U_7_land_1_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_7;
  reg FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_2_sva_2;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_2_sva_2;
  reg IsNaN_6U_10U_7_land_2_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_7;
  reg FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_3_sva_2;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_3_sva_2;
  reg IsNaN_6U_10U_7_land_3_lpi_1_dfm_3;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_7;
  reg FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_4;
  reg [3:0] FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3;
  reg [22:0] FpAdd_6U_10U_3_a_int_mant_p1_sva_2;
  reg [22:0] FpAdd_6U_10U_3_b_int_mant_p1_sva_2;
  reg IsNaN_6U_10U_7_land_lpi_1_dfm_3;
  reg [9:0] FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6;
  reg [9:0] FpAdd_6U_10U_3_o_mant_lpi_1_dfm_7;
  reg [16:0] m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2;
  reg [16:0] m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2;
  reg [16:0] m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2;
  reg [16:0] m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2;
  reg [16:0] m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2;
  reg [16:0] m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2;
  reg [16:0] m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2;
  reg [16:0] m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2;
  reg data_truncate_equal_tmp_3;
  reg data_truncate_equal_tmp_4;
  reg data_truncate_nor_tmp_4;
  reg data_truncate_nor_tmp_5;
  reg data_truncate_nor_dfs_3;
  reg data_truncate_nor_dfs_4;
  reg m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st;
  reg m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st;
  reg m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st;
  reg m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_land_lpi_1_dfm_st;
  reg m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st;
  reg m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st;
  reg m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st;
  reg m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st;
  reg m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st;
  reg m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st;
  reg m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st;
  reg m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_4_land_lpi_1_dfm_st;
  reg m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st;
  reg m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st;
  reg m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st;
  reg m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_6_land_lpi_1_dfm_st;
  reg o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm;
  reg o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2;
  reg o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st;
  reg o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm;
  reg o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2;
  reg o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_st;
  reg IsNaN_6U_10U_9_nor_1_itm;
  reg IsNaN_6U_10U_9_nor_1_itm_2;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm_2;
  reg o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm;
  reg o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2;
  reg o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_st;
  reg IsNaN_6U_10U_9_nor_2_itm;
  reg IsNaN_6U_10U_9_nor_2_itm_2;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm_2;
  reg o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm;
  reg o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2;
  reg o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_st;
  reg IsNaN_6U_10U_9_nor_3_itm;
  reg IsNaN_6U_10U_9_nor_3_itm_2;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm;
  reg IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm_2;
  reg o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st;
  reg o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st;
  reg o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st;
  reg o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st;
  reg o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm;
  reg o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_12_land_1_lpi_1_dfm_st;
  reg o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm;
  reg o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_12_land_2_lpi_1_dfm_st;
  reg IsNaN_6U_10U_13_nor_1_itm;
  reg IsNaN_6U_10U_13_nor_1_itm_2;
  reg IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm;
  reg IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2;
  reg o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm;
  reg o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_12_land_3_lpi_1_dfm_st;
  reg o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm;
  reg o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_12_land_lpi_1_dfm_st;
  reg o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm;
  reg o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm;
  reg o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2;
  reg o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_14_land_1_lpi_1_dfm_st;
  reg o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm;
  reg o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm;
  reg o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2;
  reg o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_14_land_2_lpi_1_dfm_st;
  reg o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm;
  reg o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm;
  reg o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2;
  reg o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_14_land_3_lpi_1_dfm_st;
  reg o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm;
  reg o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm;
  reg o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2;
  reg o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st;
  reg IsNaN_6U_10U_14_land_lpi_1_dfm_st;
  reg [16:0] IntSubExt_16U_16U_17U_o_acc_1_itm;
  reg [16:0] IntSubExt_16U_16U_17U_o_acc_1_itm_2;
  reg [16:0] IntAddExt_16U_16U_17U_o_acc_itm;
  reg [16:0] IntAddExt_16U_16U_17U_o_acc_itm_2;
  reg [16:0] IntSubExt_16U_16U_17U_1_o_acc_1_itm;
  reg [16:0] IntSubExt_16U_16U_17U_1_o_acc_1_itm_2;
  reg [16:0] IntSubExt_16U_16U_17U_2_o_acc_1_itm;
  reg [16:0] IntSubExt_16U_16U_17U_2_o_acc_1_itm_2;
  reg [16:0] IntSubExt_16U_16U_17U_o_acc_2_itm;
  reg [16:0] IntSubExt_16U_16U_17U_o_acc_2_itm_2;
  reg [16:0] IntAddExt_16U_16U_17U_o_acc_1_itm;
  reg [16:0] IntAddExt_16U_16U_17U_o_acc_1_itm_2;
  reg [16:0] IntSubExt_16U_16U_17U_1_o_acc_2_itm;
  reg [16:0] IntSubExt_16U_16U_17U_1_o_acc_2_itm_2;
  reg [16:0] IntSubExt_16U_16U_17U_2_o_acc_2_itm;
  reg [16:0] IntSubExt_16U_16U_17U_2_o_acc_2_itm_2;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  reg data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm;
  reg data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  reg data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg IsNaN_6U_10U_16_nor_12_itm;
  reg IsNaN_6U_10U_16_nor_12_itm_2;
  reg IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm;
  reg IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm_2;
  reg data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st;
  reg IsNaN_6U_10U_16_nor_15_itm;
  reg IsNaN_6U_10U_16_nor_15_itm_2;
  reg IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm;
  reg IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm_2;
  reg data_truncate_mux1h_410_itm_3;
  reg data_truncate_mux1h_410_itm_4;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_404_itm_3;
  reg data_truncate_mux1h_404_itm_4;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_398_itm_3;
  reg data_truncate_mux1h_398_itm_4;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_392_itm_3;
  reg data_truncate_mux1h_392_itm_4;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_386_itm_3;
  reg data_truncate_mux1h_386_itm_4;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_380_itm_3;
  reg data_truncate_mux1h_380_itm_4;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_374_itm_3;
  reg data_truncate_mux1h_374_itm_4;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_368_itm_3;
  reg data_truncate_mux1h_368_itm_4;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_362_itm_3;
  reg data_truncate_mux1h_362_itm_4;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_356_itm_3;
  reg data_truncate_mux1h_356_itm_4;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_350_itm_3;
  reg data_truncate_mux1h_350_itm_4;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_344_itm_3;
  reg data_truncate_mux1h_344_itm_4;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_338_itm_3;
  reg data_truncate_mux1h_338_itm_4;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_332_itm_3;
  reg data_truncate_mux1h_332_itm_4;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_326_itm_3;
  reg data_truncate_mux1h_326_itm_4;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg data_truncate_mux1h_320_itm_3;
  reg data_truncate_mux1h_320_itm_4;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
  reg IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
  reg data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4;
  reg data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
  reg data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_2;
  reg IsNaN_6U_10U_4_land_lpi_1_dfm_st_2;
  reg o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
  reg o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4;
  reg o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4;
  reg o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_st_4;
  reg o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
  reg o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  reg IsNaN_6U_10U_10_land_1_lpi_1_dfm_st_3;
  reg o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
  reg o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  reg IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3;
  reg o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
  reg IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3;
  reg o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
  reg o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  reg IsNaN_6U_10U_10_land_lpi_1_dfm_st_3;
  reg o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
  reg o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4;
  reg IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_4;
  reg o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_4;
  reg o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_4;
  reg o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_12_land_lpi_1_dfm_st_3;
  reg IsNaN_6U_10U_12_land_lpi_1_dfm_st_4;
  reg o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_14_land_1_lpi_1_dfm_st_4;
  reg o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_14_land_2_lpi_1_dfm_st_4;
  reg o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
  reg IsNaN_6U_10U_14_land_3_lpi_1_dfm_st_4;
  reg o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
  reg o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4;
  reg IsNaN_6U_10U_14_land_lpi_1_dfm_st_4;
  reg data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  reg FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_1;
  reg FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_0;
  reg FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_1;
  reg FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_0;
  reg FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_1;
  reg FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_0;
  reg FpAdd_6U_10U_qr_5_4_lpi_1_dfm_1;
  reg FpAdd_6U_10U_qr_5_4_lpi_1_dfm_0;
  reg FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_1;
  reg FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_0;
  reg FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_1;
  reg FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_0;
  reg FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_1;
  reg FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_0;
  reg FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_1;
  reg FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_0;
  reg FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_1;
  reg FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_0;
  reg FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_1;
  reg FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_0;
  reg FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_1;
  reg FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_0;
  reg FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_1;
  reg FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_0;
  reg FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_1;
  reg FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_0;
  reg FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_1;
  reg FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_0;
  reg FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_1;
  reg FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_0;
  reg FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_1;
  reg FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_0_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_16U_mbits_fixed_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_1_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_2_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_3_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_4_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_5_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_6_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_7_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_8_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_9_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_10_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_11_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_12_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_13_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_14_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_15_sva_1_20_2_1;
  reg [18:0] IntShiftRight_18U_2U_8U_mbits_fixed_sva_1_20_2_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_0_1;
  wire and_1769_cse;
  wire and_1771_cse;
  wire and_1801_cse;
  wire and_1803_cse;
  wire and_1833_cse;
  wire and_1835_cse;
  wire and_1865_cse;
  wire and_1867_cse;
  wire and_1895_cse;
  wire and_1897_cse;
  wire and_1927_cse;
  wire and_1929_cse;
  wire and_1959_cse;
  wire and_1961_cse;
  wire and_1991_cse;
  wire and_1993_cse;
  wire and_2021_cse;
  wire and_2023_cse;
  wire and_2053_cse;
  wire and_2055_cse;
  wire and_2085_cse;
  wire and_2087_cse;
  wire and_2117_cse;
  wire and_2119_cse;
  wire and_2147_cse;
  wire and_2149_cse;
  wire and_2179_cse;
  wire and_2181_cse;
  wire and_2211_cse;
  wire and_2213_cse;
  wire and_2243_cse;
  wire and_2245_cse;
  wire main_stage_en_1;
  wire IsDenorm_5U_10U_7_land_lpi_1_dfm;
  wire IsInf_5U_10U_7_land_lpi_1_dfm;
  wire IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_sva;
  wire IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_sva;
  wire IsDenorm_5U_10U_7_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_7_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_3_sva;
  wire IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_3_sva;
  wire IsDenorm_5U_10U_7_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_7_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_2_sva;
  wire IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_2_sva;
  wire IsDenorm_5U_10U_7_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_7_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_1_sva;
  wire IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_1_sva;
  wire IsDenorm_5U_10U_2_land_lpi_1_dfm;
  wire IsInf_5U_10U_2_land_lpi_1_dfm;
  wire IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva;
  wire IsDenorm_5U_10U_2_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_2_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_3_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva;
  wire IsDenorm_5U_10U_2_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_2_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_2_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva;
  wire IsDenorm_5U_10U_2_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_2_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_1_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva;
  wire IsDenorm_5U_10U_1_land_lpi_1_dfm;
  wire IsInf_5U_10U_1_land_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva;
  wire IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_sva;
  wire IsDenorm_5U_10U_land_lpi_1_dfm;
  wire IsInf_5U_10U_land_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva;
  wire IsDenorm_5U_10U_1_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_1_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva;
  wire IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_3_sva;
  wire IsDenorm_5U_10U_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva;
  wire IsDenorm_5U_10U_1_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_1_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva;
  wire IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_2_sva;
  wire IsDenorm_5U_10U_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva;
  wire IsDenorm_5U_10U_1_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_1_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva;
  wire IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_1_sva;
  wire IsDenorm_5U_10U_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva;
  wire FpAdd_6U_10U_3_and_25_ssc;
  wire FpAdd_6U_10U_3_and_10_tmp;
  wire FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_6_m1c;
  wire FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_3_and_23_ssc;
  wire FpAdd_6U_10U_3_and_9_tmp;
  wire FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_5_m1c;
  wire FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_3_and_21_ssc;
  wire FpAdd_6U_10U_3_and_8_tmp;
  wire FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_4_m1c;
  wire FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_2_and_25_ssc;
  wire FpAdd_6U_10U_2_and_10_tmp;
  wire FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_6_m1c;
  wire FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_2_and_23_ssc;
  wire FpAdd_6U_10U_2_and_9_tmp;
  wire FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_5_m1c;
  wire FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_2_and_21_ssc;
  wire FpAdd_6U_10U_2_and_8_tmp;
  wire FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_4_m1c;
  wire FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_1_and_25_ssc;
  wire FpAdd_6U_10U_1_and_10_tmp;
  wire FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_6_m1c;
  wire FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_1_and_23_ssc;
  wire FpAdd_6U_10U_1_and_9_tmp;
  wire FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_5_m1c;
  wire FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_1_and_21_ssc;
  wire FpAdd_6U_10U_1_and_8_tmp;
  wire FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_4_m1c;
  wire FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_and_25_ssc;
  wire FpAdd_6U_10U_and_10_tmp;
  wire FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_6_m1c;
  wire FpAdd_6U_10U_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_and_23_ssc;
  wire FpAdd_6U_10U_and_9_tmp;
  wire FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  wire FpAdd_6U_10U_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_and_21_ssc;
  wire FpAdd_6U_10U_and_8_tmp;
  wire FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_4_m1c;
  wire FpAdd_6U_10U_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_3_and_27_ssc;
  wire FpAdd_6U_10U_3_and_11_tmp;
  wire FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_7_m1c;
  wire FpAdd_6U_10U_3_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_2_and_27_ssc;
  wire FpAdd_6U_10U_2_and_11_tmp;
  wire FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_7_m1c;
  wire FpAdd_6U_10U_2_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_1_and_27_ssc;
  wire FpAdd_6U_10U_1_and_11_tmp;
  wire FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  wire FpAdd_6U_10U_1_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_and_27_ssc;
  wire FpAdd_6U_10U_and_11_tmp;
  wire FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  wire FpAdd_6U_10U_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_9_m1c;
  wire FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_7_m1c;
  wire FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_5_m1c;
  wire FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_9_m1c;
  wire FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_7_m1c;
  wire FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_5_m1c;
  wire FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_9_m1c;
  wire FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_7_m1c;
  wire FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_5_m1c;
  wire FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_9_m1c;
  wire FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_7_m1c;
  wire FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_5_m1c;
  wire FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_11_m1c;
  wire FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_11_m1c;
  wire FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_11_m1c;
  wire FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_11_m1c;
  wire FpAdd_6U_10U_7_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_6_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_5_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_4_is_inf_lpi_1_dfm;
  wire FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm;
  wire FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm;
  wire FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm;
  wire FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_o_sign_2_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_1_mx0;
  wire FpAdd_6U_10U_o_sign_3_lpi_1_dfm_1_mx0;
  wire data_truncate_equal_tmp_mx0w0;
  wire data_truncate_nor_tmp_mx0w0;
  wire FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_o_expo_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_4_mx0;
  wire FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_mx0;
  wire FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_4_mx0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1;
  wire [3:0] FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_3_int_mant_p1_sva;
  wire [3:0] FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_3_int_mant_p1_3_sva;
  wire [3:0] FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_3_int_mant_p1_2_sva;
  wire [3:0] FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_3_int_mant_p1_1_sva;
  wire [3:0] FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_2_int_mant_p1_sva;
  wire [3:0] FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_2_int_mant_p1_3_sva;
  wire [3:0] FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_2_int_mant_p1_2_sva;
  wire [3:0] FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_2_int_mant_p1_1_sva;
  wire [3:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_sva;
  wire [3:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_3_sva;
  wire [3:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_2_sva;
  wire [3:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_1_sva;
  wire [3:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_sva;
  wire [3:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_3_sva;
  wire [3:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_2_sva;
  wire [3:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_1_sva;
  wire [5:0] FpAdd_6U_10U_7_o_expo_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_6_o_expo_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_5_o_expo_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_4_o_expo_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_2;
  wire [5:0] FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_3_int_mant_p1_sva_1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_3_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_3_int_mant_p1_3_sva_1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_2_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_3_int_mant_p1_2_sva_1;
  wire [23:0] FpAdd_6U_10U_3_int_mant_p1_1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_3_int_mant_p1_1_sva_1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_2_int_mant_p1_sva_1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_3_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_2_int_mant_p1_3_sva_1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_2_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_2_int_mant_p1_2_sva_1;
  wire [23:0] FpAdd_6U_10U_2_int_mant_p1_1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_2_int_mant_p1_1_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_int_mant_p1_sva_1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_3_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_int_mant_p1_3_sva_1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_2_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_int_mant_p1_2_sva_1;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_int_mant_p1_1_sva_1;
  wire m_row0_m_row0_nor_3_m1c;
  wire m_row0_m_row0_nor_15_m1c;
  wire m_row0_m_row0_nor_14_m1c;
  wire m_row0_m_row0_nor_13_m1c;
  wire m_row0_m_row0_nor_2_m1c;
  wire m_row0_m_row0_nor_12_m1c;
  wire m_row0_m_row0_nor_11_m1c;
  wire m_row0_m_row0_nor_10_m1c;
  wire m_row0_m_row0_nor_1_m1c;
  wire m_row0_m_row0_nor_9_m1c;
  wire m_row0_m_row0_nor_8_m1c;
  wire m_row0_m_row0_nor_7_m1c;
  wire m_row0_m_row0_nor_m1c;
  wire m_row0_m_row0_nor_6_m1c;
  wire m_row0_m_row0_nor_5_m1c;
  wire m_row0_m_row0_nor_4_m1c;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_1_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_2_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_3_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_4_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_5_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_6_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_7_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_8_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_9_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_10_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_11_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_12_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_13_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_14_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_15_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_8U_mbits_fixed_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_1_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_2_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_3_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_4_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_5_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_6_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_7_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_8_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_9_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_10_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_11_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_12_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_13_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_14_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_15_tmp;
  reg [18:0] reg_IntShiftRight_18U_2U_16U_mbits_fixed_tmp;
  wire and_1474_m1c;
  wire and_1469_m1c;
  wire and_1459_m1c;
  wire and_1454_m1c;
  wire and_1449_m1c;
  wire and_1439_m1c;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2;
  wire chn_data_out_and_cse;
  wire nor_57_cse;
  wire or_181_cse;
  reg reg_chn_data_out_rsci_ld_core_psct_cse;
  wire or_317_cse;
  wire nor_150_cse;
  wire or_427_cse;
  wire or_429_cse;
  wire or_434_cse;
  wire or_476_cse;
  wire and_2507_cse;
  wire and_2491_cse;
  wire and_2495_cse;
  wire IsNaN_6U_10U_16_and_cse;
  wire IsNaN_6U_10U_12_aelse_and_cse;
  wire or_99_cse;
  wire or_109_cse;
  wire or_119_cse;
  wire or_256_cse;
  wire or_237_cse;
  wire or_209_cse;
  wire or_196_cse;
  wire or_183_cse;
  wire nor_82_cse;
  wire or_152_cse;
  wire nor_70_cse;
  wire FpAdd_6U_10U_3_b_int_mant_p1_and_cse;
  wire IsNaN_6U_10U_6_aelse_and_cse;
  wire FpAdd_6U_10U_3_and_29_cse;
  wire FpAdd_6U_10U_3_and_32_cse;
  wire FpAdd_6U_10U_3_and_35_cse;
  wire FpAdd_6U_10U_3_and_38_cse;
  wire FpAdd_6U_10U_2_and_29_cse;
  wire FpAdd_6U_10U_2_and_32_cse;
  wire FpAdd_6U_10U_2_and_35_cse;
  wire FpAdd_6U_10U_2_and_38_cse;
  wire FpAdd_6U_10U_1_and_29_cse;
  wire FpAdd_6U_10U_1_and_32_cse;
  wire FpAdd_6U_10U_1_and_35_cse;
  wire FpAdd_6U_10U_1_and_38_cse;
  wire FpAdd_6U_10U_and_29_cse;
  wire FpAdd_6U_10U_and_32_cse;
  wire FpAdd_6U_10U_and_35_cse;
  wire FpAdd_6U_10U_and_38_cse;
  wire or_623_cse;
  wire or_648_cse;
  wire or_638_cse;
  wire or_629_cse;
  wire IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse;
  wire IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_cse;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_cse;
  wire IntSubExt_16U_16U_17U_2_o_and_cse;
  wire [9:0] m_row2_if_d1_mux_1_cse;
  wire [9:0] m_row2_if_d1_mux_4_cse;
  wire [9:0] m_row2_if_d1_mux_7_cse;
  wire nor_384_cse;
  wire nor_562_cse;
  wire nor_559_cse;
  wire nor_555_cse;
  wire nor_551_cse;
  wire nor_545_cse;
  wire nor_540_cse;
  wire nor_535_cse;
  wire or_796_cse;
  wire or_311_cse;
  wire or_315_cse;
  wire and_2555_cse;
  wire and_2550_cse;
  wire and_2545_cse;
  wire or_371_cse;
  wire or_373_cse;
  wire or_375_cse;
  wire and_2537_cse;
  wire and_2532_cse;
  wire and_2527_cse;
  wire and_2517_cse;
  wire and_2512_cse;
  wire and_2503_cse;
  wire and_2498_cse;
  wire and_2487_cse;
  wire or_548_cse;
  wire and_2481_cse;
  wire or_567_cse;
  wire and_2475_cse;
  wire and_2464_cse;
  wire or_87_cse;
  wire FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1;
  wire FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1;
  wire FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1;
  wire FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1;
  wire FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1;
  wire FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1;
  wire FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1;
  wire FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1;
  wire FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1;
  wire FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1;
  wire FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1;
  wire FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1;
  wire FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1;
  wire FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1;
  wire FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1;
  wire FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1;
  wire nand_147_cse;
  wire or_527_cse;
  wire or_134_cse;
  wire and_828_cse;
  wire or_325_cse;
  wire and_2556_cse;
  wire and_72_cse;
  wire or_521_cse;
  wire or_224_cse;
  wire mux_13_cse;
  wire mux_16_cse;
  wire mux_40_cse;
  wire FpAdd_6U_10U_3_b_int_mant_p1_and_4_cse;
  wire mux_24_cse;
  wire mux_46_cse;
  wire mux_cse;
  wire mux_9_cse;
  wire mux_11_cse;
  wire mux_27_cse;
  wire mux_29_cse;
  wire mux_31_cse;
  wire mux_33_cse;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0;
  wire [20:0] IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0;
  wire and_358_rgt;
  wire and_360_rgt;
  wire and_370_rgt;
  wire and_374_rgt;
  wire and_383_rgt;
  wire and_386_rgt;
  wire and_388_rgt;
  wire and_390_rgt;
  wire and_392_rgt;
  wire and_401_rgt;
  wire and_404_rgt;
  wire and_413_rgt;
  wire and_416_rgt;
  wire and_418_rgt;
  wire and_420_rgt;
  wire and_422_rgt;
  wire and_431_rgt;
  wire and_434_rgt;
  wire and_443_rgt;
  wire and_446_rgt;
  wire and_448_rgt;
  wire and_450_rgt;
  wire and_452_rgt;
  wire and_454_rgt;
  wire and_456_rgt;
  wire and_459_rgt;
  wire and_461_rgt;
  wire and_463_rgt;
  wire and_466_rgt;
  wire and_468_rgt;
  wire and_470_rgt;
  wire and_473_rgt;
  wire and_475_rgt;
  wire and_477_rgt;
  wire and_479_rgt;
  wire and_481_rgt;
  wire and_484_rgt;
  wire and_486_rgt;
  wire and_488_rgt;
  wire and_491_rgt;
  wire and_493_rgt;
  wire and_495_rgt;
  wire and_498_rgt;
  wire and_500_rgt;
  wire and_502_rgt;
  wire and_504_rgt;
  wire and_506_rgt;
  wire and_509_rgt;
  wire and_511_rgt;
  wire and_513_rgt;
  wire and_516_rgt;
  wire and_518_rgt;
  wire and_520_rgt;
  wire and_523_rgt;
  wire and_525_rgt;
  wire and_527_rgt;
  wire and_537_rgt;
  wire and_540_rgt;
  wire and_548_rgt;
  wire and_551_rgt;
  wire and_564_rgt;
  wire and_567_rgt;
  wire and_575_rgt;
  wire and_578_rgt;
  wire and_590_rgt;
  wire and_593_rgt;
  wire and_601_rgt;
  wire and_604_rgt;
  wire and_610_rgt;
  wire and_612_rgt;
  wire and_614_rgt;
  wire and_616_rgt;
  wire and_620_rgt;
  wire and_622_rgt;
  wire and_624_rgt;
  wire and_626_rgt;
  wire and_630_rgt;
  wire and_632_rgt;
  wire and_634_rgt;
  wire and_636_rgt;
  wire and_640_rgt;
  wire and_642_rgt;
  wire and_644_rgt;
  wire and_646_rgt;
  wire and_649_rgt;
  wire and_652_rgt;
  wire and_654_rgt;
  wire and_656_rgt;
  wire and_658_rgt;
  wire and_661_rgt;
  wire and_664_rgt;
  wire and_666_rgt;
  wire and_668_rgt;
  wire and_670_rgt;
  wire and_673_rgt;
  wire and_676_rgt;
  wire and_680_rgt;
  wire and_683_rgt;
  wire and_689_rgt;
  wire and_691_rgt;
  wire and_693_rgt;
  wire and_695_rgt;
  wire and_697_rgt;
  wire and_699_rgt;
  wire and_701_rgt;
  wire and_703_rgt;
  wire and_705_rgt;
  wire and_707_rgt;
  wire and_709_rgt;
  wire and_711_rgt;
  wire and_713_rgt;
  wire and_715_rgt;
  wire and_717_rgt;
  wire and_719_rgt;
  wire and_721_rgt;
  wire and_723_rgt;
  wire and_725_rgt;
  wire and_727_rgt;
  wire and_733_rgt;
  wire and_735_rgt;
  wire and_737_rgt;
  wire and_739_rgt;
  wire and_741_rgt;
  wire and_743_rgt;
  wire and_745_rgt;
  wire and_747_rgt;
  wire and_749_rgt;
  wire and_751_rgt;
  wire and_753_rgt;
  wire and_755_rgt;
  wire and_757_rgt;
  wire and_759_rgt;
  wire and_761_rgt;
  wire and_763_rgt;
  wire and_765_rgt;
  wire and_767_rgt;
  wire and_769_rgt;
  wire and_771_rgt;
  wire and_773_rgt;
  wire and_775_rgt;
  wire and_777_rgt;
  wire and_779_rgt;
  wire and_781_rgt;
  wire and_783_rgt;
  wire and_785_rgt;
  wire and_787_rgt;
  wire and_789_rgt;
  wire and_791_rgt;
  wire and_793_rgt;
  wire and_795_rgt;
  wire and_932_rgt;
  wire and_935_rgt;
  wire and_938_rgt;
  wire and_941_rgt;
  wire and_946_rgt;
  wire and_949_rgt;
  wire and_952_rgt;
  wire and_955_rgt;
  wire and_960_rgt;
  wire and_963_rgt;
  wire and_966_rgt;
  wire and_969_rgt;
  wire and_974_rgt;
  wire and_977_rgt;
  wire and_980_rgt;
  wire and_983_rgt;
  wire and_985_rgt;
  wire and_988_rgt;
  wire and_991_rgt;
  wire and_994_rgt;
  wire and_997_rgt;
  wire and_999_rgt;
  wire and_1002_rgt;
  wire and_1005_rgt;
  wire and_1008_rgt;
  wire and_1011_rgt;
  wire and_1013_rgt;
  wire and_1016_rgt;
  wire and_1019_rgt;
  wire and_1022_rgt;
  wire and_1025_rgt;
  wire and_1030_rgt;
  wire and_1033_rgt;
  wire and_1036_rgt;
  wire and_1039_rgt;
  wire and_1044_rgt;
  wire and_1047_rgt;
  wire and_1050_rgt;
  wire and_1053_rgt;
  wire and_1058_rgt;
  wire and_1061_rgt;
  wire and_1064_rgt;
  wire and_1067_rgt;
  wire and_1069_rgt;
  wire and_1072_rgt;
  wire and_1075_rgt;
  wire and_1078_rgt;
  wire and_1081_rgt;
  wire and_1083_rgt;
  wire and_1086_rgt;
  wire and_1089_rgt;
  wire and_1092_rgt;
  wire and_1095_rgt;
  wire and_1097_rgt;
  wire and_1268_rgt;
  wire and_1271_rgt;
  wire and_1280_rgt;
  wire and_1283_rgt;
  wire and_1285_rgt;
  wire and_1288_rgt;
  wire and_1291_rgt;
  wire and_1294_rgt;
  wire and_1303_rgt;
  wire and_1306_rgt;
  wire and_1314_rgt;
  wire and_1317_rgt;
  wire and_1323_rgt;
  wire and_1325_rgt;
  wire and_1327_rgt;
  wire and_1329_rgt;
  wire and_1333_rgt;
  wire and_1335_rgt;
  wire and_1337_rgt;
  wire and_1339_rgt;
  wire and_1342_rgt;
  wire and_1345_rgt;
  wire and_1348_rgt;
  wire and_1351_rgt;
  wire and_1354_rgt;
  wire and_1357_rgt;
  wire and_1362_rgt;
  wire and_1365_rgt;
  wire and_1368_rgt;
  wire and_1371_rgt;
  wire and_1373_rgt;
  wire and_1376_rgt;
  wire and_1379_rgt;
  wire and_1382_rgt;
  wire and_1385_rgt;
  wire and_1390_rgt;
  wire and_1393_rgt;
  wire and_1396_rgt;
  wire and_1399_rgt;
  wire and_1401_rgt;
  wire FpAdd_6U_10U_o_sign_or_1_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_1_rgt;
  wire m_row1_if_d2_or_1_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_4_rgt;
  wire FpAdd_6U_10U_o_sign_or_11_rgt;
  wire and_1440_rgt;
  wire and_1442_rgt;
  wire and_1444_rgt;
  wire m_row1_if_d2_or_11_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_17_rgt;
  wire FpAdd_6U_10U_o_sign_or_8_rgt;
  wire and_1460_rgt;
  wire and_1462_rgt;
  wire and_1464_rgt;
  wire m_row1_if_d2_or_8_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_14_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_9_rgt;
  wire m_row1_if_d2_or_3_rgt;
  wire FpAdd_6U_10U_1_o_sign_or_6_rgt;
  wire FpAdd_6U_10U_o_sign_or_3_rgt;
  wire [9:0] m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm;
  wire [9:0] m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm;
  wire [9:0] m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm;
  wire [9:0] m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm;
  wire [9:0] m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm;
  wire [9:0] m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm;
  wire [9:0] m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm;
  wire [9:0] m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm;
  wire [22:0] m_row0_1_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] m_row0_2_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] m_row0_3_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] m_row0_4_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] m_row1_1_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [22:0] m_row1_2_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [22:0] m_row1_3_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [22:0] m_row1_4_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [22:0] m_row2_1_FpNormalize_6U_23U_2_else_lshift_itm;
  wire [22:0] m_row2_2_FpNormalize_6U_23U_2_else_lshift_itm;
  wire [22:0] m_row2_3_FpNormalize_6U_23U_2_else_lshift_itm;
  wire [22:0] m_row2_4_FpNormalize_6U_23U_2_else_lshift_itm;
  wire [22:0] m_row3_1_FpNormalize_6U_23U_3_else_lshift_itm;
  wire [22:0] m_row3_2_FpNormalize_6U_23U_3_else_lshift_itm;
  wire [22:0] m_row3_3_FpNormalize_6U_23U_3_else_lshift_itm;
  wire [22:0] m_row3_4_FpNormalize_6U_23U_3_else_lshift_itm;
  wire [22:0] o_col0_1_FpNormalize_6U_23U_4_else_lshift_itm;
  wire [22:0] o_col0_2_FpNormalize_6U_23U_4_else_lshift_itm;
  wire [22:0] o_col0_3_FpNormalize_6U_23U_4_else_lshift_itm;
  wire [22:0] o_col0_4_FpNormalize_6U_23U_4_else_lshift_itm;
  wire [22:0] o_col1_1_FpNormalize_6U_23U_5_else_lshift_itm;
  wire [22:0] o_col1_2_FpNormalize_6U_23U_5_else_lshift_itm;
  wire [22:0] o_col1_3_FpNormalize_6U_23U_5_else_lshift_itm;
  wire [22:0] o_col1_4_FpNormalize_6U_23U_5_else_lshift_itm;
  wire [22:0] o_col2_1_FpNormalize_6U_23U_6_else_lshift_itm;
  wire [22:0] o_col2_2_FpNormalize_6U_23U_6_else_lshift_itm;
  wire [22:0] o_col2_3_FpNormalize_6U_23U_6_else_lshift_itm;
  wire [22:0] o_col2_4_FpNormalize_6U_23U_6_else_lshift_itm;
  wire [22:0] o_col3_1_FpNormalize_6U_23U_7_else_lshift_itm;
  wire [22:0] o_col3_2_FpNormalize_6U_23U_7_else_lshift_itm;
  wire [22:0] o_col3_3_FpNormalize_6U_23U_7_else_lshift_itm;
  wire [22:0] o_col3_4_FpNormalize_6U_23U_7_else_lshift_itm;
  wire [10:0] data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire [10:0] data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm;
  wire FpAdd_6U_10U_mux_3_itm;
  wire FpAdd_6U_10U_mux_20_itm;
  wire FpAdd_6U_10U_mux_37_itm;
  wire FpAdd_6U_10U_mux_69_itm;
  wire FpAdd_6U_10U_1_mux_3_itm;
  wire FpAdd_6U_10U_1_mux_20_itm;
  wire FpAdd_6U_10U_1_mux_37_itm;
  wire FpAdd_6U_10U_1_mux_73_itm;
  wire FpAdd_6U_10U_2_mux_3_itm;
  wire FpAdd_6U_10U_2_mux_20_itm;
  wire FpAdd_6U_10U_2_mux_37_itm;
  wire FpAdd_6U_10U_2_mux_73_itm;
  wire FpAdd_6U_10U_3_mux_3_itm;
  wire FpAdd_6U_10U_3_mux_20_itm;
  wire FpAdd_6U_10U_3_mux_37_itm;
  wire FpAdd_6U_10U_3_mux_69_itm;
  wire [17:0] z_out;
  wire [18:0] nl_z_out;
  wire [17:0] z_out_1;
  wire [18:0] nl_z_out_1;
  wire [17:0] z_out_2;
  wire [18:0] nl_z_out_2;
  wire [17:0] z_out_3;
  wire [18:0] nl_z_out_3;
  wire [17:0] z_out_4;
  wire [18:0] nl_z_out_4;
  wire [17:0] z_out_5;
  wire [18:0] nl_z_out_5;
  wire [17:0] z_out_6;
  wire [18:0] nl_z_out_6;
  wire [17:0] z_out_7;
  wire [18:0] nl_z_out_7;
  wire [17:0] z_out_8;
  wire [18:0] nl_z_out_8;
  wire [17:0] z_out_9;
  wire [18:0] nl_z_out_9;
  wire [17:0] z_out_10;
  wire [18:0] nl_z_out_10;
  wire [17:0] z_out_11;
  wire [18:0] nl_z_out_11;
  wire [17:0] z_out_12;
  wire [18:0] nl_z_out_12;
  wire [17:0] z_out_13;
  wire [18:0] nl_z_out_13;
  wire [17:0] z_out_14;
  wire [18:0] nl_z_out_14;
  wire [17:0] z_out_15;
  wire [18:0] nl_z_out_15;
  wire FpAdd_6U_10U_7_if_2_and_tmp;
  wire FpAdd_6U_10U_7_if_2_and_tmp_1;
  wire FpAdd_6U_10U_7_if_2_and_tmp_2;
  wire FpAdd_6U_10U_7_if_2_and_tmp_3;
  wire FpAdd_6U_10U_6_if_2_and_tmp;
  wire FpAdd_6U_10U_6_if_2_and_tmp_1;
  wire FpAdd_6U_10U_6_if_2_and_tmp_2;
  wire FpAdd_6U_10U_6_if_2_and_tmp_3;
  wire FpAdd_6U_10U_5_if_2_and_tmp;
  wire FpAdd_6U_10U_5_if_2_and_tmp_1;
  wire FpAdd_6U_10U_5_if_2_and_tmp_2;
  wire FpAdd_6U_10U_5_if_2_and_tmp_3;
  wire FpAdd_6U_10U_4_if_2_and_tmp;
  wire FpAdd_6U_10U_4_if_2_and_tmp_1;
  wire FpAdd_6U_10U_4_if_2_and_tmp_2;
  wire FpAdd_6U_10U_4_if_2_and_tmp_3;
  wire chn_data_in_rsci_ld_core_psct_mx0c0;
  wire m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  wire o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  wire data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  wire main_stage_v_1_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w4;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_2_mx0w4;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w4;
  wire m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_a_int_mant_p1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_b_int_mant_p1_sva_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_4_mx0w4;
  wire m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_a_int_mant_p1_3_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_b_int_mant_p1_3_sva_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_2_mx0w4;
  wire m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_a_int_mant_p1_2_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_b_int_mant_p1_2_sva_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_mx0w4;
  wire m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_a_int_mant_p1_1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_3_b_int_mant_p1_1_sva_mx0w0;
  wire m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_a_int_mant_p1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_b_int_mant_p1_sva_mx0w0;
  wire m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_a_int_mant_p1_3_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_b_int_mant_p1_3_sva_mx0w0;
  wire m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_a_int_mant_p1_2_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_b_int_mant_p1_2_sva_mx0w0;
  wire m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_a_int_mant_p1_1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_2_b_int_mant_p1_1_sva_mx0w0;
  wire m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_a_int_mant_p1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_b_int_mant_p1_sva_mx0w0;
  wire m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_a_int_mant_p1_3_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_b_int_mant_p1_3_sva_mx0w0;
  wire m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_a_int_mant_p1_2_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_b_int_mant_p1_2_sva_mx0w0;
  wire m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_a_int_mant_p1_1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_1_b_int_mant_p1_1_sva_mx0w0;
  wire m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_a_int_mant_p1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_b_int_mant_p1_sva_mx0w0;
  wire m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_a_int_mant_p1_3_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_b_int_mant_p1_3_sva_mx0w0;
  wire m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_a_int_mant_p1_2_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_b_int_mant_p1_2_sva_mx0w0;
  wire m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
  wire [22:0] FpAdd_6U_10U_a_int_mant_p1_1_sva_mx0w0;
  wire [22:0] FpAdd_6U_10U_b_int_mant_p1_1_sva_mx0w0;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire [9:0] FpAdd_6U_10U_7_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_7_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_7_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_6_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_6_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_6_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_5_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_5_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_5_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_4_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_4_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpAdd_6U_10U_4_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_8_mx0w0;
  wire [5:0] FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_7_o_mant_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_7_o_expo_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_6_o_mant_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_6_o_expo_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_5_o_mant_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_5_o_expo_lpi_1_dfm_8_mx0w0;
  wire [9:0] FpAdd_6U_10U_4_o_mant_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpAdd_6U_10U_4_o_expo_lpi_1_dfm_8_mx0w0;
  wire FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx0c1;
  wire [9:0] FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx1;
  wire FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx0c1;
  wire [9:0] FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx1;
  wire FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx0c1;
  wire [9:0] FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx1;
  wire FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0c1;
  wire [9:0] FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_3_mx0;
  wire FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_qr_3_0_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_mx0c1;
  wire FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_6_mx0w4;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_6_mx0w4;
  wire o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
  wire o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
  wire o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
  wire o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
  wire o_col1_4_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
  wire o_col1_3_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
  wire o_col1_2_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
  wire o_col1_1_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
  wire o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
  wire o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
  wire o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
  wire o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
  wire o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
  wire o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
  wire o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
  wire o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
  wire data_truncate_nor_dfs_mx0w0;
  wire IsNaN_6U_10U_9_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_9_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_9_land_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0;
  wire [1:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_3_mx0;
  wire o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
  wire o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
  wire o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
  wire o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
  wire o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
  wire o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
  wire o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
  wire o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
  wire o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
  wire o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
  wire o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
  wire o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
  wire o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
  wire o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
  wire o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
  wire o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
  wire FpAdd_6U_10U_4_mux_45_mx1w1;
  wire FpAdd_6U_10U_4_mux_13_mx1w1;
  wire FpAdd_6U_10U_5_mux_45_mx1w1;
  wire FpAdd_6U_10U_5_mux_13_mx1w1;
  wire FpAdd_6U_10U_6_mux_45_mx1w1;
  wire FpAdd_6U_10U_6_mux_13_mx1w1;
  wire FpAdd_6U_10U_4_mux_29_mx1w1;
  wire FpAdd_6U_10U_5_mux_29_mx1w1;
  wire FpAdd_6U_10U_6_mux_29_mx1w1;
  wire FpAdd_6U_10U_4_mux_61_mx1w1;
  wire FpAdd_6U_10U_5_mux_61_mx1w1;
  wire FpAdd_6U_10U_6_mux_61_mx1w1;
  wire data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
  wire FpAdd_6U_10U_7_mux_13_mx1w0;
  wire FpAdd_6U_10U_7_mux_29_mx1w0;
  wire FpAdd_6U_10U_7_mux_45_mx1w0;
  wire FpAdd_6U_10U_7_mux_61_mx1w0;
  wire FpAdd_6U_10U_o_sign_1_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_1_mux_19_mx0w2;
  wire FpAdd_6U_10U_1_mux_36_mx0w2;
  wire FpAdd_6U_10U_3_o_sign_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_2_o_sign_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_1_o_sign_lpi_1_dfm_3_mx0c2;
  wire FpAdd_6U_10U_o_sign_lpi_1_dfm_3_mx0c2;
  wire [16:0] IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0;
  wire [16:0] m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
  wire [16:0] IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0;
  wire [16:0] m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
  wire [16:0] IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0;
  wire [18:0] nl_IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0;
  wire [16:0] m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [16:0] IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0;
  wire [16:0] m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [16:0] m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
  wire [16:0] m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
  wire [16:0] m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [16:0] m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [17:0] nl_m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
  wire [16:0] IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0;
  wire [16:0] IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0;
  wire [16:0] IntAddExt_16U_16U_17U_o_acc_itm_mx0w0;
  wire [18:0] nl_IntAddExt_16U_16U_17U_o_acc_itm_mx0w0;
  wire [16:0] IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0;
  wire [17:0] nl_IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_3_cse;
  wire IsNaN_5U_10U_7_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_cse;
  wire IsNaN_5U_10U_2_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_2_cse;
  wire IsNaN_5U_10U_7_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_cse;
  wire IsNaN_5U_10U_2_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_1_cse;
  wire IsNaN_5U_10U_7_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_cse;
  wire IsNaN_5U_10U_2_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_cse;
  wire IsNaN_5U_10U_7_land_1_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_cse;
  wire IsNaN_5U_10U_2_land_1_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse;
  wire IsNaN_5U_10U_1_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse;
  wire IsNaN_5U_10U_1_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse;
  wire IsNaN_5U_10U_1_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse;
  wire IsNaN_5U_10U_1_land_1_lpi_1_dfm;
  wire IsZero_5U_10U_2_land_lpi_1_dfm;
  wire IsZero_5U_10U_2_land_3_lpi_1_dfm;
  wire IsZero_5U_10U_2_land_2_lpi_1_dfm;
  wire IsZero_5U_10U_2_land_1_lpi_1_dfm;
  wire IsZero_5U_10U_1_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse;
  wire IsNaN_5U_10U_land_lpi_1_dfm;
  wire IsZero_5U_10U_1_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse;
  wire IsNaN_5U_10U_land_3_lpi_1_dfm;
  wire IsZero_5U_10U_1_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse;
  wire IsNaN_5U_10U_land_2_lpi_1_dfm;
  wire IsZero_5U_10U_1_land_1_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse;
  wire IsNaN_5U_10U_land_1_lpi_1_dfm;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_1_sva;
  wire [5:0] FpAdd_6U_10U_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_1_sva_4;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_2_sva;
  wire [5:0] FpAdd_6U_10U_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_2_sva_4;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_3_sva;
  wire [5:0] FpAdd_6U_10U_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_3_sva_4;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_1_else_carry_1_sva;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_1_sva_4;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_1_else_carry_2_sva;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_2_sva_4;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_1_else_carry_3_sva;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_3_sva_4;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_1_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_2_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_2_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_2_else_carry_1_sva;
  wire [5:0] FpAdd_6U_10U_2_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_1_sva_4;
  wire [22:0] FpAdd_6U_10U_2_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_2_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_2_else_carry_2_sva;
  wire [5:0] FpAdd_6U_10U_2_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_2_sva_4;
  wire [22:0] FpAdd_6U_10U_2_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_2_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_2_else_carry_3_sva;
  wire [5:0] FpAdd_6U_10U_2_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_3_sva_4;
  wire [22:0] FpAdd_6U_10U_2_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_2_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_2_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_2_o_expo_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_3_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_3_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_3_else_carry_1_sva;
  wire [5:0] FpAdd_6U_10U_3_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_1_sva_4;
  wire [22:0] FpAdd_6U_10U_3_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_3_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_3_else_carry_2_sva;
  wire [5:0] FpAdd_6U_10U_3_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_2_sva_4;
  wire [22:0] FpAdd_6U_10U_3_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_3_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [21:0] FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_3_else_carry_3_sva;
  wire [5:0] FpAdd_6U_10U_3_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_3_sva_4;
  wire [22:0] FpAdd_6U_10U_3_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_3_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_3_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_3_o_expo_lpi_1_dfm_1;
  wire [9:0] FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_2_mx0;
  wire [9:0] FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0;
  wire [9:0] FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5;
  wire FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_4;
  wire [3:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0;
  wire FpMantRNE_23U_11U_3_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpAdd_6U_10U_3_and_24_ssc;
  wire FpAdd_6U_10U_3_and_17_ssc;
  wire FpAdd_6U_10U_3_and_22_ssc;
  wire FpAdd_6U_10U_3_and_15_ssc;
  wire FpAdd_6U_10U_3_and_20_ssc;
  wire FpAdd_6U_10U_3_and_13_ssc;
  wire FpMantRNE_23U_11U_2_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpAdd_6U_10U_2_and_24_ssc;
  wire FpAdd_6U_10U_2_and_17_ssc;
  wire FpAdd_6U_10U_2_and_22_ssc;
  wire FpAdd_6U_10U_2_and_15_ssc;
  wire FpAdd_6U_10U_2_and_20_ssc;
  wire FpAdd_6U_10U_2_and_13_ssc;
  wire FpMantRNE_23U_11U_1_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpAdd_6U_10U_1_and_24_ssc;
  wire FpAdd_6U_10U_1_and_17_ssc;
  wire FpAdd_6U_10U_1_and_22_ssc;
  wire FpAdd_6U_10U_1_and_15_ssc;
  wire FpAdd_6U_10U_1_and_20_ssc;
  wire FpAdd_6U_10U_1_and_13_ssc;
  wire FpMantRNE_23U_11U_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpAdd_6U_10U_and_24_ssc;
  wire FpAdd_6U_10U_and_17_ssc;
  wire FpAdd_6U_10U_and_22_ssc;
  wire FpAdd_6U_10U_and_15_ssc;
  wire FpAdd_6U_10U_and_20_ssc;
  wire FpAdd_6U_10U_and_13_ssc;
  wire [22:0] FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_1;
  wire [22:0] FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_1;
  wire FpMantRNE_23U_11U_7_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_7_else_carry_3_sva;
  wire [21:0] FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_7_else_carry_2_sva;
  wire [21:0] FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_7_else_carry_1_sva;
  wire [21:0] FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_6_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_6_else_carry_3_sva;
  wire [21:0] FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_6_else_carry_2_sva;
  wire [21:0] FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_6_else_carry_1_sva;
  wire [21:0] FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_5_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_5_else_carry_3_sva;
  wire [21:0] FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_5_else_carry_2_sva;
  wire [21:0] FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_5_else_carry_1_sva;
  wire [21:0] FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_4_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_4_else_carry_3_sva;
  wire [21:0] FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_4_else_carry_2_sva;
  wire [21:0] FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_4_else_carry_1_sva;
  wire [21:0] FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire IsNaN_6U_10U_16_land_lpi_1_dfm;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_3_mx0;
  wire IsNaN_6U_10U_16_land_13_lpi_1_dfm;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_1_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_1_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_1_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_1_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_1_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_2_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_2_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_2_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_2_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_2_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_3_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_3_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_3_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_3_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_3_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_4_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_4_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_4_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_4_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_4_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_5_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_5_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_5_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_5_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_5_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_6_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_6_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_6_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_6_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_6_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_7_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_7_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_7_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_7_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_7_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_8_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_8_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_8_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_8_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_8_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_9_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_9_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_9_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_9_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_9_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_10_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_10_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_10_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_10_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_10_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_11_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_11_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_11_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_11_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_11_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_12_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_12_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_12_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_12_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_12_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_13_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_13_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_13_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_13_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_13_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_14_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_14_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_14_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_14_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_14_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_15_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_15_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_15_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_15_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_15_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva;
  wire [2:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva;
  wire [3:0] nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_guard_mask_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_stick_mask_sva;
  wire [11:0] nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_sva;
  wire [9:0] FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_sva;
  wire [10:0] FpMantDecShiftRight_10U_6U_10U_least_mask_sva;
  wire FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_5;
  wire [3:0] FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_3_0;
  wire FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_4;
  wire FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_5;
  wire [3:0] FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_3_0;
  wire FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_4;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5;
  wire [3:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4;
  wire FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5;
  wire [3:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0;
  wire FpAdd_6U_10U_o_expo_lpi_1_dfm_7_4;
  wire [5:0] FpAdd_6U_10U_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_sva_4;
  wire [5:0] FpAdd_6U_10U_1_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_sva_4;
  wire [5:0] FpAdd_6U_10U_2_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_2_o_expo_sva_4;
  wire [5:0] FpAdd_6U_10U_3_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_3_o_expo_sva_4;
  wire FpAdd_6U_10U_3_and_26_ssc;
  wire FpAdd_6U_10U_3_and_19_ssc;
  wire FpAdd_6U_10U_2_and_26_ssc;
  wire FpAdd_6U_10U_2_and_19_ssc;
  wire FpAdd_6U_10U_1_and_26_ssc;
  wire FpAdd_6U_10U_1_and_19_ssc;
  wire FpAdd_6U_10U_and_26_ssc;
  wire FpAdd_6U_10U_and_19_ssc;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_asn_19_mx0w1;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_a_int_mant_p1_1_sva;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_asn_13_mx0w1;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_a_int_mant_p1_2_sva;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_asn_7_mx0w1;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_a_int_mant_p1_3_sva;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_asn_1_mx0w1;
  wire [22:0] FpAdd_6U_10U_4_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_4_a_int_mant_p1_sva;
  wire [5:0] FpAdd_6U_10U_5_b_right_shift_qr_1_sva;
  wire [7:0] nl_FpAdd_6U_10U_5_b_right_shift_qr_1_sva;
  wire [5:0] FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1;
  wire [7:0] nl_FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_asn_19_mx0w1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_a_int_mant_p1_1_sva;
  wire [5:0] FpAdd_6U_10U_5_b_right_shift_qr_2_sva;
  wire [7:0] nl_FpAdd_6U_10U_5_b_right_shift_qr_2_sva;
  wire [5:0] FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1;
  wire [7:0] nl_FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_asn_13_mx0w1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_a_int_mant_p1_2_sva;
  wire [5:0] FpAdd_6U_10U_5_b_right_shift_qr_3_sva;
  wire [7:0] nl_FpAdd_6U_10U_5_b_right_shift_qr_3_sva;
  wire [5:0] FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1;
  wire [7:0] nl_FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_asn_7_mx0w1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_a_int_mant_p1_3_sva;
  wire [5:0] FpAdd_6U_10U_5_b_right_shift_qr_sva;
  wire [7:0] nl_FpAdd_6U_10U_5_b_right_shift_qr_sva;
  wire [5:0] FpAdd_6U_10U_5_a_right_shift_qr_sva_1;
  wire [7:0] nl_FpAdd_6U_10U_5_a_right_shift_qr_sva_1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_asn_1_mx0w1;
  wire [22:0] FpAdd_6U_10U_5_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_5_a_int_mant_p1_sva;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_asn_19_mx0w1;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_a_int_mant_p1_1_sva;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_asn_13_mx0w1;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_a_int_mant_p1_2_sva;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_asn_7_mx0w1;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_a_int_mant_p1_3_sva;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_asn_1_mx0w1;
  wire [22:0] FpAdd_6U_10U_6_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_6_a_int_mant_p1_sva;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_asn_19_mx0w1;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_a_int_mant_p1_1_sva;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_asn_13_mx0w1;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_a_int_mant_p1_2_sva;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_asn_7_mx0w1;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_a_int_mant_p1_3_sva;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_asn_1_mx0w1;
  wire [22:0] FpAdd_6U_10U_7_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_7_a_int_mant_p1_sva;
  wire FpAdd_6U_10U_7_and_3_tmp;
  wire FpAdd_6U_10U_7_and_2_tmp;
  wire FpAdd_6U_10U_7_and_1_tmp;
  wire FpAdd_6U_10U_7_and_tmp;
  wire FpAdd_6U_10U_6_and_3_tmp;
  wire FpAdd_6U_10U_6_and_2_tmp;
  wire FpAdd_6U_10U_6_and_1_tmp;
  wire FpAdd_6U_10U_6_and_tmp;
  wire FpAdd_6U_10U_5_and_3_tmp;
  wire FpAdd_6U_10U_5_and_2_tmp;
  wire FpAdd_6U_10U_5_and_1_tmp;
  wire FpAdd_6U_10U_5_and_tmp;
  wire FpAdd_6U_10U_4_and_3_tmp;
  wire FpAdd_6U_10U_4_and_2_tmp;
  wire FpAdd_6U_10U_4_and_1_tmp;
  wire FpAdd_6U_10U_4_and_tmp;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_15_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_15_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_14_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_14_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_13_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_13_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_12_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_12_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_11_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_11_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_10_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_10_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_9_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_9_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_8_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_8_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_7_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_7_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_6_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_6_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_5_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_5_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_4_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_4_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_3_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_3_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_2_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_2_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_1_sva;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_1_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_19;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_19;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_21;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_21;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_23;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_23;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_25;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_25;
  wire m_row1_1_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2;
  wire m_row1_2_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2;
  wire m_row1_3_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2;
  wire m_row1_4_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2;
  wire m_row2_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2;
  wire m_row2_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2;
  wire m_row2_3_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2;
  wire m_row2_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2;
  wire IsZero_5U_10U_7_aelse_not_13;
  wire IsZero_5U_10U_7_aelse_not_15;
  wire IsZero_5U_10U_7_aelse_not_17;
  wire IsZero_5U_10U_7_aelse_not_19;
  wire IsZero_5U_10U_aelse_not_13;
  wire IsZero_5U_10U_aelse_not_15;
  wire IsZero_5U_10U_aelse_not_17;
  wire IsZero_5U_10U_aelse_not_19;
  wire m_row2_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2;
  wire m_row2_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2;
  wire m_row2_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2;
  wire m_row2_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2;
  wire FpNormalize_6U_23U_oelse_not_9;
  wire FpNormalize_6U_23U_oelse_not_11;
  wire FpNormalize_6U_23U_oelse_not_13;
  wire FpNormalize_6U_23U_oelse_not_15;
  wire FpNormalize_6U_23U_1_oelse_not_9;
  wire FpNormalize_6U_23U_1_oelse_not_11;
  wire FpNormalize_6U_23U_1_oelse_not_13;
  wire FpNormalize_6U_23U_1_oelse_not_15;
  wire FpNormalize_6U_23U_2_oelse_not_9;
  wire FpNormalize_6U_23U_2_oelse_not_11;
  wire FpNormalize_6U_23U_2_oelse_not_13;
  wire FpNormalize_6U_23U_2_oelse_not_15;
  wire FpNormalize_6U_23U_3_oelse_not_9;
  wire FpNormalize_6U_23U_3_oelse_not_11;
  wire FpNormalize_6U_23U_3_oelse_not_13;
  wire FpNormalize_6U_23U_3_oelse_not_15;
  wire FpNormalize_6U_23U_4_oelse_not_9;
  wire FpNormalize_6U_23U_4_oelse_not_11;
  wire FpNormalize_6U_23U_4_oelse_not_13;
  wire FpNormalize_6U_23U_4_oelse_not_15;
  wire FpNormalize_6U_23U_5_oelse_not_9;
  wire FpNormalize_6U_23U_5_oelse_not_11;
  wire FpNormalize_6U_23U_5_oelse_not_13;
  wire FpNormalize_6U_23U_5_oelse_not_15;
  wire FpNormalize_6U_23U_6_oelse_not_9;
  wire FpNormalize_6U_23U_6_oelse_not_11;
  wire FpNormalize_6U_23U_6_oelse_not_13;
  wire FpNormalize_6U_23U_6_oelse_not_15;
  wire FpNormalize_6U_23U_7_oelse_not_9;
  wire FpNormalize_6U_23U_7_oelse_not_11;
  wire FpNormalize_6U_23U_7_oelse_not_13;
  wire FpNormalize_6U_23U_7_oelse_not_15;
  wire m_row0_asn_184;
  wire m_row0_asn_186;
  wire m_row0_asn_188;
  wire m_row0_asn_190;
  wire m_row0_asn_192;
  wire m_row0_asn_194;
  wire m_row0_asn_196;
  wire m_row0_asn_198;
  wire m_row0_asn_200;
  wire m_row0_asn_202;
  wire m_row0_asn_204;
  wire m_row0_asn_206;
  wire m_row0_asn_208;
  wire m_row0_asn_210;
  wire m_row0_asn_212;
  wire m_row0_asn_214;
  wire m_row0_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2;
  wire m_row0_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2;
  wire m_row0_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2;
  wire m_row0_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2;
  wire [22:0] FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0;
  wire [22:0] FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0;
  wire m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10;
  wire m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10;
  wire m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10;
  wire m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10;
  wire m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10;
  wire m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10;
  wire m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10;
  wire m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_32;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_33;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_34;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_35;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_36;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_37;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_38;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_39;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_40;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_41;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_42;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_43;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_44;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_45;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_46;
  wire [3:0] libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_47;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_32;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_33;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_34;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_35;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_36;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_37;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_38;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_39;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_40;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_41;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_42;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_43;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_44;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_45;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_46;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_47;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_48;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_49;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_50;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_51;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_52;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_53;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_54;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_55;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_56;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_57;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_58;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_59;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_60;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_61;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_62;
  wire [4:0] libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_63;
  reg reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp;
  reg reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2;
  reg reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1;
  reg reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1;
  wire FpAdd_6U_10U_3_o_expo_and_13_ssc;
  reg reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2;
  reg reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_3_o_expo_and_12_ssc;
  reg reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_3_o_expo_and_11_ssc;
  reg reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_o_expo_and_13_ssc;
  reg reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2;
  reg reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_1_o_expo_and_13_ssc;
  reg reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2;
  reg reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_2_o_expo_and_13_ssc;
  reg reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2;
  reg reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_o_expo_and_12_ssc;
  reg reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_1_o_expo_and_12_ssc;
  reg reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_2_o_expo_and_12_ssc;
  reg reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_o_expo_and_11_ssc;
  reg reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_1_o_expo_and_11_ssc;
  reg reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_2_o_expo_and_11_ssc;
  reg reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp;
  reg reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_2;
  wire FpAdd_6U_10U_6_and_38_ssc;
  reg reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_5_and_38_ssc;
  reg reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_4_and_38_ssc;
  reg reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_6_and_42_ssc;
  reg reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_5_and_42_ssc;
  reg reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_4_and_42_ssc;
  reg reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_7_and_38_ssc;
  reg reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_7_and_42_ssc;
  reg reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_6_and_35_ssc;
  reg reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_5_and_35_ssc;
  reg reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_4_and_35_ssc;
  reg reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_6_and_39_ssc;
  reg reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_5_and_39_ssc;
  reg reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_4_and_39_ssc;
  reg reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_6_and_36_ssc;
  reg reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_5_and_36_ssc;
  reg reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_4_and_36_ssc;
  reg reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_6_and_40_ssc;
  reg reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_5_and_40_ssc;
  reg reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_4_and_40_ssc;
  reg reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_6_and_37_ssc;
  reg reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_5_and_37_ssc;
  reg reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_4_and_37_ssc;
  reg reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_6_and_41_ssc;
  reg reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_5_and_41_ssc;
  reg reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_4_and_41_ssc;
  reg reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_7_and_35_ssc;
  reg reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_7_and_39_ssc;
  reg reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_7_and_36_ssc;
  reg reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_7_and_40_ssc;
  reg reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_7_and_37_ssc;
  reg reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp;
  reg reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_2;
  wire FpAdd_6U_10U_7_and_41_ssc;
  reg reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp;
  reg reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1;
  reg [3:0] reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2;
  wire FpAdd_6U_10U_and_cse;
  wire IsNaN_6U_10U_6_aelse_and_8_cse;
  wire IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_6_cse;
  wire FpAdd_6U_10U_o_expo_and_cse;
  wire IsNaN_6U_10U_14_aelse_and_cse;
  wire IsNaN_6U_10U_16_and_4_cse;
  wire IsNaN_6U_10U_16_IsNaN_6U_10U_16_or_3_cse;
  wire FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_cse;
  wire data_truncate_and_cse;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_16_cse;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_16_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_9_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_11_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_4_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_12_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_14_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_16_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_11_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_10_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_9_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_18_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_18_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_15_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse;
  wire o_data_data_and_64_cse;
  wire o_data_data_and_80_cse;
  wire data_truncate_and_129_cse;
  wire data_truncate_and_130_cse;
  wire data_truncate_and_124_cse;
  wire data_truncate_and_125_cse;
  wire data_truncate_data_truncate_nor_1_cse;
  wire FpAdd_6U_10U_2_o_mant_and_8_cse;
  wire FpAdd_6U_10U_1_o_mant_and_8_cse;
  wire FpAdd_6U_10U_o_mant_and_8_cse;
  wire FpAdd_6U_10U_3_o_mant_and_8_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_18_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_22_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_21_cse;
  wire FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse;
  wire IntShiftRight_18U_2U_16U_mbits_fixed_and_cse;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_80_cse;
  wire IntShiftRight_18U_2U_8U_mbits_fixed_and_cse;
  wire IntShiftRight_18U_2U_8U_obits_fixed_and_144_cse;
  wire IsNaN_6U_10U_9_and_11_cse;
  wire IsNaN_6U_10U_9_and_13_cse;
  wire IsNaN_6U_10U_9_and_15_cse;
  wire IsNaN_6U_10U_13_and_3_cse;
  wire IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse;
  reg reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse;
  wire FpAdd_6U_10U_3_a_int_mant_p1_and_cse;
  wire FpAdd_6U_10U_3_a_int_mant_p1_and_7_cse;
  wire FpAdd_6U_10U_1_a_int_mant_p1_and_8_cse;
  wire IsNaN_6U_10U_12_aelse_and_4_cse;
  wire FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_16_cse;
  wire IsNaN_6U_10U_9_and_cse;
  wire IsNaN_6U_10U_9_and_7_cse;
  wire IsNaN_6U_10U_9_and_9_cse;
  wire IsNaN_6U_10U_13_and_cse;
  reg reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse;
  reg reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse;
  reg reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse;
  reg reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse;
  reg reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse;
  reg reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse;
  reg reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse;
  reg reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse;
  reg reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse;
  reg reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse;
  reg reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse;
  reg reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse;
  reg reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse;
  reg reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse;
  reg reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse;
  reg reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse;
  reg reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse;
  reg reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse;
  wire nor_439_cse;
  wire nor_546_cse;
  reg reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  reg reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  reg reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  reg reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  reg reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse;
  reg reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  reg reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  reg reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  reg reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  reg reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  reg reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  wire or_1963_cse;
  wire or_1960_cse;
  wire or_1962_cse;
  wire or_1959_cse;
  wire or_1961_cse;
  wire or_1958_cse;
  wire mux_79_cse;
  wire mux_67_cse;
  wire and_2591_cse;
  wire and_2588_cse;
  wire and_2585_cse;
  wire and_2582_cse;
  wire and_2579_cse;
  wire and_2576_cse;
  wire mux_468_cse;
  reg reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse;
  reg reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse;
  reg reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse;
  reg reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse;
  reg reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse;
  reg reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse;
  reg reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1;
  reg reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1;
  wire [9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_4_itm;
  wire [9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_5_itm;
  wire [9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_6_itm;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_4_itm;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_5_itm;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_6_itm;
  wire [9:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_4_itm;
  wire [9:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_5_itm;
  wire [9:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_6_itm;
  wire [9:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_4_itm;
  wire [9:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_5_itm;
  wire [9:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_6_itm;
  wire [9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_11_itm;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_11_itm;
  wire [9:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_11_itm;
  wire [9:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_11_itm;
  wire data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
  wire data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  wire data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  wire m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1;
  wire m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1;
  wire m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1;
  wire m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1;
  wire m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1;
  wire m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1;
  wire m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1;
  wire m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1;
  wire m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1;
  wire m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1;
  wire m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1;
  wire m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1;
  wire m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1;
  wire m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1;
  wire m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1;
  wire m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1;
  wire m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1;
  wire m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1;
  wire m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1;
  wire m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1;
  wire m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1;
  wire m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1;
  wire m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1;
  wire m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1;
  wire FpAdd_6U_10U_7_is_a_greater_acc_3_itm_6_1;
  wire FpAdd_6U_10U_7_is_a_greater_acc_2_itm_6_1;
  wire FpAdd_6U_10U_7_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_7_is_a_greater_acc_itm_6_1;
  wire FpAdd_6U_10U_6_is_a_greater_acc_3_itm_6_1;
  wire FpAdd_6U_10U_6_is_a_greater_acc_2_itm_6_1;
  wire FpAdd_6U_10U_6_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_6_is_a_greater_acc_itm_6_1;
  wire FpAdd_6U_10U_5_is_a_greater_acc_3_itm_6_1;
  wire FpAdd_6U_10U_5_is_a_greater_acc_2_itm_6_1;
  wire FpAdd_6U_10U_5_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_5_is_a_greater_acc_itm_6_1;
  wire FpAdd_6U_10U_4_is_a_greater_acc_3_itm_6_1;
  wire FpAdd_6U_10U_4_is_a_greater_acc_2_itm_6_1;
  wire FpAdd_6U_10U_4_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_4_is_a_greater_acc_itm_6_1;
  wire o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1;
  wire o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1;
  wire o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1;
  wire o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1;
  wire o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1;
  wire o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1;
  wire o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1;
  wire o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1;
  wire o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1;
  wire o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1;
  wire o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1;
  wire o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1;
  wire o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1;
  wire o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1;
  wire o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1;
  wire o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1;
  wire o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1;
  wire o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1;
  wire o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1;
  wire o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1;
  wire o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1;
  wire o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1;
  wire o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1;
  wire o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1;
  wire o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1;
  wire o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1;
  wire o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1;
  wire o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1;
  wire o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1;
  wire o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1;
  wire o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1;
  wire o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1;
  wire FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_itm_10_1;
  wire FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_itm_10_1;
  wire FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_itm_10_1;
  wire FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_itm_10_1;
  wire FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_itm_10_1;
  wire FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_itm_10_1;
  wire FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_itm_10_1;
  wire FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_itm_10_1;
  wire FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_itm_10_1;
  wire FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_itm_10_1;
  wire FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_itm_10_1;
  wire FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_itm_10_1;
  wire FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_itm_10_1;
  wire FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_itm_10_1;
  wire FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_itm_10_1;
  wire FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_itm_10_1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse;

  wire[0:0] shift_0_prb;
  wire[0:0] and_16;
  wire[0:0] shift_0_prb_1;
  wire[0:0] and_19;
  wire[0:0] shift_0_prb_2;
  wire[0:0] and_22;
  wire[0:0] shift_0_prb_3;
  wire[0:0] and_25;
  wire[0:0] shift_0_prb_4;
  wire[0:0] and_28;
  wire[0:0] shift_0_prb_5;
  wire[0:0] and_31;
  wire[0:0] shift_0_prb_6;
  wire[0:0] and_34;
  wire[0:0] shift_0_prb_7;
  wire[0:0] and_37;
  wire[0:0] shift_0_prb_8;
  wire[0:0] and_40;
  wire[0:0] shift_0_prb_9;
  wire[0:0] and_43;
  wire[0:0] shift_0_prb_10;
  wire[0:0] and_46;
  wire[0:0] shift_0_prb_11;
  wire[0:0] and_49;
  wire[0:0] shift_0_prb_12;
  wire[0:0] and_52;
  wire[0:0] shift_0_prb_13;
  wire[0:0] and_55;
  wire[0:0] shift_0_prb_14;
  wire[0:0] and_58;
  wire[0:0] shift_0_prb_15;
  wire[0:0] and_61;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_2;
  wire[0:0] iExpoWidth_oExpoWidth_prb_3;
  wire[0:0] iExpoWidth_oExpoWidth_prb_4;
  wire[0:0] iExpoWidth_oExpoWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_6;
  wire[0:0] iExpoWidth_oExpoWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_8;
  wire[0:0] iExpoWidth_oExpoWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_10;
  wire[0:0] iExpoWidth_oExpoWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_12;
  wire[0:0] iExpoWidth_oExpoWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_14;
  wire[0:0] iExpoWidth_oExpoWidth_prb_15;
  wire[0:0] iExpoWidth_oExpoWidth_prb_16;
  wire[0:0] iExpoWidth_oExpoWidth_prb_17;
  wire[0:0] iExpoWidth_oExpoWidth_prb_18;
  wire[0:0] iExpoWidth_oExpoWidth_prb_19;
  wire[0:0] iExpoWidth_oExpoWidth_prb_20;
  wire[0:0] iExpoWidth_oExpoWidth_prb_21;
  wire[0:0] iExpoWidth_oExpoWidth_prb_22;
  wire[0:0] iExpoWidth_oExpoWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_24;
  wire[0:0] iExpoWidth_oExpoWidth_prb_25;
  wire[0:0] iExpoWidth_oExpoWidth_prb_26;
  wire[0:0] iExpoWidth_oExpoWidth_prb_27;
  wire[0:0] iExpoWidth_oExpoWidth_prb_28;
  wire[0:0] iExpoWidth_oExpoWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_30;
  wire[0:0] iExpoWidth_oExpoWidth_prb_31;
  wire[0:0] oWidth_mWidth_prb;
  wire[0:0] oWidth_mWidth_prb_1;
  wire[0:0] oWidth_mWidth_prb_2;
  wire[0:0] oWidth_mWidth_prb_3;
  wire[0:0] oWidth_mWidth_prb_4;
  wire[0:0] oWidth_mWidth_prb_5;
  wire[0:0] oWidth_mWidth_prb_6;
  wire[0:0] oWidth_mWidth_prb_7;
  wire[0:0] oWidth_mWidth_prb_8;
  wire[0:0] oWidth_mWidth_prb_9;
  wire[0:0] oWidth_mWidth_prb_10;
  wire[0:0] oWidth_mWidth_prb_11;
  wire[0:0] oWidth_mWidth_prb_12;
  wire[0:0] oWidth_mWidth_prb_13;
  wire[0:0] oWidth_mWidth_prb_14;
  wire[0:0] oWidth_mWidth_prb_15;
  wire[0:0] oWidth_mWidth_prb_16;
  wire[0:0] oWidth_mWidth_prb_17;
  wire[0:0] oWidth_mWidth_prb_18;
  wire[0:0] oWidth_mWidth_prb_19;
  wire[0:0] oWidth_mWidth_prb_20;
  wire[0:0] oWidth_mWidth_prb_21;
  wire[0:0] oWidth_mWidth_prb_22;
  wire[0:0] oWidth_mWidth_prb_23;
  wire[0:0] oWidth_mWidth_prb_24;
  wire[0:0] oWidth_mWidth_prb_25;
  wire[0:0] oWidth_mWidth_prb_26;
  wire[0:0] oWidth_mWidth_prb_27;
  wire[0:0] oWidth_mWidth_prb_28;
  wire[0:0] oWidth_mWidth_prb_29;
  wire[0:0] oWidth_mWidth_prb_30;
  wire[0:0] oWidth_mWidth_prb_31;
  wire[0:0] iExpoWidth_oExpoWidth_prb_32;
  wire[0:0] iExpoWidth_oExpoWidth_prb_33;
  wire[0:0] iExpoWidth_oExpoWidth_prb_34;
  wire[0:0] iExpoWidth_oExpoWidth_prb_35;
  wire[0:0] iExpoWidth_oExpoWidth_prb_36;
  wire[0:0] iExpoWidth_oExpoWidth_prb_37;
  wire[0:0] iExpoWidth_oExpoWidth_prb_38;
  wire[0:0] iExpoWidth_oExpoWidth_prb_39;
  wire[0:0] iExpoWidth_oExpoWidth_prb_40;
  wire[0:0] iExpoWidth_oExpoWidth_prb_41;
  wire[0:0] iExpoWidth_oExpoWidth_prb_42;
  wire[0:0] iExpoWidth_oExpoWidth_prb_43;
  wire[0:0] iExpoWidth_oExpoWidth_prb_44;
  wire[0:0] iExpoWidth_oExpoWidth_prb_45;
  wire[0:0] iExpoWidth_oExpoWidth_prb_46;
  wire[0:0] iExpoWidth_oExpoWidth_prb_47;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_1_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_172_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_2_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_6_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_255_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_1_nl;
  wire[0:0] or_1299_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_1_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_3_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_17_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_5_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_17_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_256_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_2_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_3_nl;
  wire[0:0] or_1305_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_3_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_5_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_28_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_8_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_28_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_257_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_4_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_5_nl;
  wire[0:0] or_1311_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_5_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_7_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_39_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_11_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_39_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_258_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_6_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_7_nl;
  wire[0:0] or_1317_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_7_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_9_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_50_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_14_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_50_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_259_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_8_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_9_nl;
  wire[0:0] or_1323_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_9_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_11_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_61_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_17_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_61_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_260_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_10_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_11_nl;
  wire[0:0] or_1329_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_11_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_13_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_72_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_20_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_72_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_261_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_12_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_13_nl;
  wire[0:0] or_1335_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_13_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_15_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_83_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_23_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_83_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_262_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_14_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_15_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_15_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_17_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_94_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_26_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_94_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_263_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_16_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_17_nl;
  wire[0:0] or_1347_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_17_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_19_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_105_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_29_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_105_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_264_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_18_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_19_nl;
  wire[0:0] or_1353_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_19_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_21_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_116_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_32_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_116_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_265_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_20_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_21_nl;
  wire[0:0] or_1359_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_21_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_23_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_127_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_35_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_127_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_266_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_22_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_23_nl;
  wire[0:0] or_1365_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_23_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_25_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_138_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_38_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_138_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_267_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_24_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_25_nl;
  wire[0:0] or_1371_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_25_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_27_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_149_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_41_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_149_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_268_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_26_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_27_nl;
  wire[0:0] or_1377_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_27_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_29_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_160_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_44_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_160_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_269_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_28_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_29_nl;
  wire[0:0] or_1383_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_29_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_31_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_mux_171_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_47_nl;
  wire[3:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_171_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_270_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_30_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_31_nl;
  wire[0:0] or_1389_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_31_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] or_170_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] and_85_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] and_88_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] and_91_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] and_96_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] and_99_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] or_1980_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] and_100_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_13_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_13_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_13_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_13_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_11_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_11_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_11_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_11_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_10_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_10_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_10_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_10_nl;
  wire[24:0] acc_16_nl;
  wire[25:0] nl_acc_16_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_8_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_9_nl;
  wire[24:0] acc_17_nl;
  wire[25:0] nl_acc_17_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_10_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_11_nl;
  wire[24:0] acc_18_nl;
  wire[25:0] nl_acc_18_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_12_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_13_nl;
  wire[24:0] acc_19_nl;
  wire[25:0] nl_acc_19_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_14_nl;
  wire[22:0] FpAdd_6U_10U_7_else_2_mux_15_nl;
  wire[24:0] acc_20_nl;
  wire[25:0] nl_acc_20_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_8_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_9_nl;
  wire[24:0] acc_21_nl;
  wire[25:0] nl_acc_21_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_10_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_11_nl;
  wire[24:0] acc_22_nl;
  wire[25:0] nl_acc_22_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_12_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_13_nl;
  wire[24:0] acc_23_nl;
  wire[25:0] nl_acc_23_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_14_nl;
  wire[22:0] FpAdd_6U_10U_6_else_2_mux_15_nl;
  wire[24:0] acc_24_nl;
  wire[25:0] nl_acc_24_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_8_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_9_nl;
  wire[24:0] acc_25_nl;
  wire[25:0] nl_acc_25_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_10_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_11_nl;
  wire[24:0] acc_26_nl;
  wire[25:0] nl_acc_26_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_12_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_13_nl;
  wire[24:0] acc_27_nl;
  wire[25:0] nl_acc_27_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_14_nl;
  wire[22:0] FpAdd_6U_10U_5_else_2_mux_15_nl;
  wire[24:0] acc_28_nl;
  wire[25:0] nl_acc_28_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_8_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_9_nl;
  wire[24:0] acc_29_nl;
  wire[25:0] nl_acc_29_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_10_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_11_nl;
  wire[24:0] acc_30_nl;
  wire[25:0] nl_acc_30_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_12_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_13_nl;
  wire[24:0] acc_31_nl;
  wire[25:0] nl_acc_31_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_14_nl;
  wire[22:0] FpAdd_6U_10U_4_else_2_mux_15_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] and_2625_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] and_2567_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] and_2562_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] and_2561_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] or_316_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] or_319_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] or_327_nl;
  wire[0:0] or_330_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] or_331_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] or_336_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] or_344_nl;
  wire[0:0] or_347_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] or_348_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] or_353_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] or_361_nl;
  wire[0:0] or_364_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] or_365_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] and_2543_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] and_2542_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] and_2541_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] or_376_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] or_384_nl;
  wire[0:0] or_387_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] or_388_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] or_393_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] or_401_nl;
  wire[0:0] or_404_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] or_405_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] or_410_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] or_418_nl;
  wire[0:0] or_421_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] or_422_nl;
  wire[0:0] nand_46_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] and_2525_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] or_433_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] or_436_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] or_444_nl;
  wire[0:0] or_447_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] or_448_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] or_458_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] or_466_nl;
  wire[0:0] or_469_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] or_470_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_475_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] or_478_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] or_481_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] or_482_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] or_490_nl;
  wire[0:0] or_493_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] or_494_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] or_502_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] or_510_nl;
  wire[0:0] or_513_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] or_514_nl;
  wire[0:0] nand_50_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] or_522_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] or_525_nl;
  wire[0:0] or_523_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] or_529_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] or_530_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] or_538_nl;
  wire[0:0] or_541_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] or_542_nl;
  wire[0:0] nand_52_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] and_2485_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] or_549_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] or_557_nl;
  wire[0:0] or_560_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] or_561_nl;
  wire[0:0] nand_53_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] and_2479_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] or_568_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] or_576_nl;
  wire[0:0] or_579_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] or_580_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] or_588_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] or_591_nl;
  wire[0:0] or_589_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] or_595_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] or_596_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] or_604_nl;
  wire[0:0] or_607_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] or_608_nl;
  wire[0:0] nand_56_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_8_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_8_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_8_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_nl;
  wire[0:0] nand_nl;
  wire[0:0] and_2619_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_3_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_15_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] or_14_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] and_2618_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] and_2616_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nand_9_nl;
  wire[0:0] and_2615_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] and_2462_nl;
  wire[0:0] nand_133_nl;
  wire[0:0] or_613_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] and_2614_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nand_13_nl;
  wire[0:0] and_2613_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] and_2461_nl;
  wire[0:0] nand_132_nl;
  wire[0:0] or_615_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] and_2612_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] and_2460_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] and_2609_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] and_2608_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] and_2607_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] or_48_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] and_2605_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] and_2604_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] or_52_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_56_nl;
  wire[0:0] and_74_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] or_60_nl;
  wire[0:0] and_75_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] nand_150_nl;
  wire[0:0] or_62_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] or_617_nl;
  wire[0:0] and_125_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] and_2459_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] and_126_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] and_2632_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] and_127_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] and_2633_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] nor_593_nl;
  wire[5:0] data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] nor_446_nl;
  wire[5:0] data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[5:0] data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl;
  wire[3:0] data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl;
  wire[2:0] data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] and_2638_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] and_2624_nl;
  wire[0:0] or_738_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] and_2622_nl;
  wire[0:0] or_753_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] and_2620_nl;
  wire[0:0] or_768_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] or_795_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] or_840_nl;
  wire[0:0] or_847_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] or_856_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] or_855_nl;
  wire[0:0] or_857_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] or_861_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] or_871_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] or_870_nl;
  wire[0:0] or_872_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] or_917_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] or_916_nl;
  wire[0:0] or_918_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_355_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] nor_351_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] and_2617_nl;
  wire[0:0] nand_19_nl;
  wire[0:0] and_2611_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] nand_21_nl;
  wire[0:0] and_2610_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] and_2425_nl;
  wire[0:0] nand_123_nl;
  wire[0:0] or_942_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] and_2606_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] and_2603_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] and_2602_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] or_69_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] nand_71_nl;
  wire[0:0] and_2424_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] or_944_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] or_945_nl;
  wire[0:0] or_946_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] or_948_nl;
  wire[0:0] or_951_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] or_953_nl;
  wire[0:0] or_954_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] or_956_nl;
  wire[0:0] or_959_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] or_961_nl;
  wire[0:0] or_962_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] or_964_nl;
  wire[0:0] or_967_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] or_970_nl;
  wire[0:0] or_971_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] or_974_nl;
  wire[0:0] or_975_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] or_978_nl;
  wire[0:0] or_979_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] or_985_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] or_986_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] and_2423_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_349_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] and_2422_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] nor_348_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] and_2421_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] nor_347_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] nor_346_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] or_999_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] or_1000_nl;
  wire[0:0] or_998_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] or_1003_nl;
  wire[0:0] or_1004_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] or_1006_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] nand_77_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] nor_345_nl;
  wire[0:0] nand_118_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] nand_116_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] nor_342_nl;
  wire[0:0] nand_115_nl;
  wire[0:0] and_337_nl;
  wire[0:0] and_339_nl;
  wire[0:0] or_1110_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_33_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_18_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_37_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_3_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_16_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_24_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_31_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_6_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_14_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_25_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl;
  wire[10:0] FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_3_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_3_is_a_greater_acc_3_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_31_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_6_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_14_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_25_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_6_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_8_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_22_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_8_nl;
  wire[10:0] FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_3_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_3_is_a_greater_acc_2_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_35_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_3_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_16_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_24_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_5_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_24_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_5_nl;
  wire[10:0] FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_3_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_3_is_a_greater_acc_1_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_37_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_18_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_26_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_2_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_26_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_2_nl;
  wire[10:0] FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl;
  wire[6:0] FpAdd_6U_10U_3_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_3_is_a_greater_acc_nl;
  wire[10:0] FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_2_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_2_is_a_greater_acc_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_8_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_8_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_22_nl;
  wire[10:0] FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_2_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_2_is_a_greater_acc_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_6_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_5_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_24_nl;
  wire[10:0] FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_2_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_2_is_a_greater_acc_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_4_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_2_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_26_nl;
  wire[10:0] FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl;
  wire[6:0] FpAdd_6U_10U_2_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_2_is_a_greater_acc_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_nl;
  wire[6:0] data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl;
  wire[5:0] data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl;
  wire[6:0] data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[6:0] data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[7:0] nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl;
  wire[9:0] FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_10_nl;
  wire[9:0] o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[10:0] nl_o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[0:0] m_row0_and_49_nl;
  wire[0:0] m_row0_and_50_nl;
  wire[9:0] FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_9_nl;
  wire[9:0] o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[10:0] nl_o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[0:0] m_row0_and_51_nl;
  wire[0:0] m_row0_and_52_nl;
  wire[9:0] FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_8_nl;
  wire[9:0] o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[10:0] nl_o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[0:0] m_row0_and_53_nl;
  wire[0:0] m_row0_and_54_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[6:0] nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_31_nl;
  wire[0:0] FpAdd_6U_10U_7_and_19_nl;
  wire[0:0] FpAdd_6U_10U_7_and_32_nl;
  wire[0:0] FpAdd_6U_10U_7_and_21_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[6:0] nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_29_nl;
  wire[0:0] FpAdd_6U_10U_7_and_13_nl;
  wire[0:0] FpAdd_6U_10U_7_and_30_nl;
  wire[0:0] FpAdd_6U_10U_7_and_15_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[6:0] nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_nl;
  wire[0:0] FpAdd_6U_10U_7_and_6_nl;
  wire[0:0] FpAdd_6U_10U_7_and_28_nl;
  wire[0:0] FpAdd_6U_10U_7_and_9_nl;
  wire[9:0] FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_10_nl;
  wire[9:0] o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[10:0] nl_o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[0:0] m_row0_and_57_nl;
  wire[0:0] m_row0_and_58_nl;
  wire[9:0] FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_9_nl;
  wire[9:0] o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[10:0] nl_o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[0:0] m_row0_and_59_nl;
  wire[0:0] m_row0_and_60_nl;
  wire[9:0] FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_8_nl;
  wire[9:0] o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[10:0] nl_o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[0:0] m_row0_and_61_nl;
  wire[0:0] m_row0_and_62_nl;
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[6:0] nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_31_nl;
  wire[0:0] FpAdd_6U_10U_6_and_19_nl;
  wire[0:0] FpAdd_6U_10U_6_and_32_nl;
  wire[0:0] FpAdd_6U_10U_6_and_21_nl;
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[6:0] nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_29_nl;
  wire[0:0] FpAdd_6U_10U_6_and_13_nl;
  wire[0:0] FpAdd_6U_10U_6_and_30_nl;
  wire[0:0] FpAdd_6U_10U_6_and_15_nl;
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[6:0] nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_nl;
  wire[0:0] FpAdd_6U_10U_6_and_6_nl;
  wire[0:0] FpAdd_6U_10U_6_and_28_nl;
  wire[0:0] FpAdd_6U_10U_6_and_9_nl;
  wire[9:0] FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_10_nl;
  wire[9:0] o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[10:0] nl_o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[0:0] m_row0_and_65_nl;
  wire[0:0] m_row0_and_66_nl;
  wire[9:0] FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_9_nl;
  wire[9:0] o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[10:0] nl_o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[0:0] m_row0_and_67_nl;
  wire[0:0] m_row0_and_68_nl;
  wire[9:0] FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_8_nl;
  wire[9:0] o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[10:0] nl_o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[0:0] m_row0_and_69_nl;
  wire[0:0] m_row0_and_70_nl;
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[6:0] nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_31_nl;
  wire[0:0] FpAdd_6U_10U_5_and_19_nl;
  wire[0:0] FpAdd_6U_10U_5_and_32_nl;
  wire[0:0] FpAdd_6U_10U_5_and_21_nl;
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[6:0] nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_29_nl;
  wire[0:0] FpAdd_6U_10U_5_and_13_nl;
  wire[0:0] FpAdd_6U_10U_5_and_30_nl;
  wire[0:0] FpAdd_6U_10U_5_and_15_nl;
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[6:0] nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_nl;
  wire[0:0] FpAdd_6U_10U_5_and_6_nl;
  wire[0:0] FpAdd_6U_10U_5_and_28_nl;
  wire[0:0] FpAdd_6U_10U_5_and_9_nl;
  wire[9:0] FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_10_nl;
  wire[9:0] o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[10:0] nl_o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[0:0] m_row0_and_73_nl;
  wire[0:0] m_row0_and_74_nl;
  wire[9:0] FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_9_nl;
  wire[9:0] o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[10:0] nl_o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[0:0] m_row0_and_75_nl;
  wire[0:0] m_row0_and_76_nl;
  wire[9:0] FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_8_nl;
  wire[9:0] o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[10:0] nl_o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[0:0] m_row0_and_77_nl;
  wire[0:0] m_row0_and_78_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[6:0] nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_31_nl;
  wire[0:0] FpAdd_6U_10U_4_and_19_nl;
  wire[0:0] FpAdd_6U_10U_4_and_32_nl;
  wire[0:0] FpAdd_6U_10U_4_and_21_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[6:0] nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_29_nl;
  wire[0:0] FpAdd_6U_10U_4_and_13_nl;
  wire[0:0] FpAdd_6U_10U_4_and_30_nl;
  wire[0:0] FpAdd_6U_10U_4_and_15_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[6:0] nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_nl;
  wire[0:0] FpAdd_6U_10U_4_and_6_nl;
  wire[0:0] FpAdd_6U_10U_4_and_28_nl;
  wire[0:0] FpAdd_6U_10U_4_and_9_nl;
  wire[9:0] FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_11_nl;
  wire[9:0] o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[10:0] nl_o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl;
  wire[0:0] m_row0_and_47_nl;
  wire[0:0] m_row0_and_48_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[6:0] nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_33_nl;
  wire[0:0] FpAdd_6U_10U_7_and_25_nl;
  wire[0:0] FpAdd_6U_10U_7_and_34_nl;
  wire[0:0] FpAdd_6U_10U_7_and_27_nl;
  wire[9:0] FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_11_nl;
  wire[9:0] o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[10:0] nl_o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl;
  wire[0:0] m_row0_and_55_nl;
  wire[0:0] m_row0_and_56_nl;
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[6:0] nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_33_nl;
  wire[0:0] FpAdd_6U_10U_6_and_25_nl;
  wire[0:0] FpAdd_6U_10U_6_and_34_nl;
  wire[0:0] FpAdd_6U_10U_6_and_27_nl;
  wire[9:0] FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_11_nl;
  wire[9:0] o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[10:0] nl_o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl;
  wire[0:0] m_row0_and_63_nl;
  wire[0:0] m_row0_and_64_nl;
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[6:0] nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_33_nl;
  wire[0:0] FpAdd_6U_10U_5_and_25_nl;
  wire[0:0] FpAdd_6U_10U_5_and_34_nl;
  wire[0:0] FpAdd_6U_10U_5_and_27_nl;
  wire[9:0] FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_11_nl;
  wire[9:0] o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[10:0] nl_o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl;
  wire[0:0] m_row0_and_71_nl;
  wire[0:0] m_row0_and_72_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[6:0] nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_33_nl;
  wire[0:0] FpAdd_6U_10U_4_and_25_nl;
  wire[0:0] FpAdd_6U_10U_4_and_34_nl;
  wire[0:0] FpAdd_6U_10U_4_and_27_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_15_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_14_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_13_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_15_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_7_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_14_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_13_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_35_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_9_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_12_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_26_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_33_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_9_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_12_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_27_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_9_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_11_nl;
  wire[0:0] IsZero_5U_10U_2_aelse_not_20_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_11_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_10_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_11_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_20_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_17_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_12_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_mux1h_8_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_or_4_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_and_3_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_mux1h_20_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_2_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_and_3_nl;
  wire[0:0] m_row1_if_d2_mux1h_4_nl;
  wire[0:0] m_row1_if_d2_or_4_nl;
  wire[0:0] m_row1_if_d2_and_3_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_mux1h_24_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_10_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_and_7_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_mux1h_11_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_or_5_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_and_7_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_mux1h_23_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_7_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_and_11_nl;
  wire[0:0] m_row1_if_d2_mux1h_7_nl;
  wire[0:0] m_row1_if_d2_or_5_nl;
  wire[0:0] m_row1_if_d2_and_7_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_mux1h_27_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_11_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_and_15_nl;
  wire[0:0] FpAdd_6U_10U_4_else_6_mux_6_nl;
  wire[0:0] FpAdd_6U_10U_4_mux_33_nl;
  wire[0:0] FpAdd_6U_10U_4_else_6_mux_nl;
  wire[0:0] FpAdd_6U_10U_4_mux_1_nl;
  wire[0:0] FpAdd_6U_10U_5_else_6_mux_6_nl;
  wire[0:0] FpAdd_6U_10U_5_mux_33_nl;
  wire[0:0] FpAdd_6U_10U_5_else_6_mux_nl;
  wire[0:0] FpAdd_6U_10U_5_mux_1_nl;
  wire[0:0] FpAdd_6U_10U_6_else_6_mux_6_nl;
  wire[0:0] FpAdd_6U_10U_6_mux_33_nl;
  wire[0:0] FpAdd_6U_10U_6_else_6_mux_nl;
  wire[0:0] FpAdd_6U_10U_6_mux_1_nl;
  wire[0:0] FpAdd_6U_10U_4_else_6_mux_3_nl;
  wire[0:0] FpAdd_6U_10U_4_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_5_else_6_mux_3_nl;
  wire[0:0] FpAdd_6U_10U_5_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_6_else_6_mux_3_nl;
  wire[0:0] FpAdd_6U_10U_6_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_4_else_6_mux_9_nl;
  wire[0:0] FpAdd_6U_10U_4_mux_49_nl;
  wire[0:0] FpAdd_6U_10U_5_else_6_mux_9_nl;
  wire[0:0] FpAdd_6U_10U_5_mux_49_nl;
  wire[0:0] FpAdd_6U_10U_6_else_6_mux_9_nl;
  wire[0:0] FpAdd_6U_10U_6_mux_49_nl;
  wire[0:0] FpAdd_6U_10U_7_else_6_mux_nl;
  wire[0:0] FpAdd_6U_10U_7_mux_1_nl;
  wire[0:0] FpAdd_6U_10U_7_else_6_mux_3_nl;
  wire[0:0] FpAdd_6U_10U_7_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_7_else_6_mux_6_nl;
  wire[0:0] FpAdd_6U_10U_7_mux_33_nl;
  wire[0:0] FpAdd_6U_10U_7_else_6_mux_9_nl;
  wire[0:0] FpAdd_6U_10U_7_mux_49_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_11_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_and_7_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_13_nl;
  wire[5:0] m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[5:0] m_row0_1_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_m_row0_1_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl;
  wire[5:0] m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] m_row0_1_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_m_row0_1_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_1_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_and_5_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_19_nl;
  wire[5:0] m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[5:0] m_row0_2_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_m_row0_2_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl;
  wire[5:0] m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] m_row0_2_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_m_row0_2_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_23_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_2_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_and_3_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_25_nl;
  wire[5:0] m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[5:0] m_row0_3_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_m_row0_3_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl;
  wire[5:0] m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] m_row0_3_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_m_row0_3_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_29_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_3_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_and_1_nl;
  wire[0:0] FpAdd_6U_10U_o_expo_mux_31_nl;
  wire[5:0] m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[5:0] m_row0_4_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_m_row0_4_FpNormalize_6U_23U_else_acc_nl;
  wire[5:0] m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_11_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_and_7_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_13_nl;
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] m_row1_1_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_m_row1_1_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl;
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[9:0] m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_1_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_and_5_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_19_nl;
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] m_row1_2_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_m_row1_2_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl;
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[9:0] m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_23_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_2_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_and_3_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_25_nl;
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] m_row1_3_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_m_row1_3_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl;
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[9:0] m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_29_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_3_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_and_1_nl;
  wire[0:0] FpAdd_6U_10U_1_o_expo_mux_31_nl;
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] m_row1_4_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_m_row1_4_FpNormalize_6U_23U_1_else_acc_nl;
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_11_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_and_7_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_13_nl;
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[5:0] m_row2_1_FpNormalize_6U_23U_2_else_acc_nl;
  wire[7:0] nl_m_row2_1_FpNormalize_6U_23U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_nl;
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[9:0] m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[10:0] nl_m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_1_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_and_5_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_19_nl;
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[5:0] m_row2_2_FpNormalize_6U_23U_2_else_acc_nl;
  wire[7:0] nl_m_row2_2_FpNormalize_6U_23U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_1_nl;
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[9:0] m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[10:0] nl_m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_23_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_2_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_and_3_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_25_nl;
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[5:0] m_row2_3_FpNormalize_6U_23U_2_else_acc_nl;
  wire[7:0] nl_m_row2_3_FpNormalize_6U_23U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_2_nl;
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[9:0] m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[10:0] nl_m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_29_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_3_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_and_1_nl;
  wire[0:0] FpAdd_6U_10U_2_o_expo_mux_31_nl;
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl;
  wire[5:0] m_row2_4_FpNormalize_6U_23U_2_else_acc_nl;
  wire[7:0] nl_m_row2_4_FpNormalize_6U_23U_2_else_acc_nl;
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_11_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_and_7_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_13_nl;
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[5:0] m_row3_1_FpNormalize_6U_23U_3_else_acc_nl;
  wire[7:0] nl_m_row3_1_FpNormalize_6U_23U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_nl;
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[9:0] m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[10:0] nl_m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_17_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_1_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_and_5_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_19_nl;
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[5:0] m_row3_2_FpNormalize_6U_23U_3_else_acc_nl;
  wire[7:0] nl_m_row3_2_FpNormalize_6U_23U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_1_nl;
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[9:0] m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[10:0] nl_m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_23_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_2_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_and_3_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_25_nl;
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[5:0] m_row3_3_FpNormalize_6U_23U_3_else_acc_nl;
  wire[7:0] nl_m_row3_3_FpNormalize_6U_23U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_2_nl;
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[9:0] m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[10:0] nl_m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_29_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_3_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_and_1_nl;
  wire[0:0] FpAdd_6U_10U_3_o_expo_mux_31_nl;
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[6:0] nl_m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl;
  wire[5:0] m_row3_4_FpNormalize_6U_23U_3_else_acc_nl;
  wire[7:0] nl_m_row3_4_FpNormalize_6U_23U_3_else_acc_nl;
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[6:0] nl_m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_13_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_2_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_13_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_2_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_13_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_2_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_11_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_1_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_11_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_1_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_1_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_11_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_1_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_9_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_9_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_9_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_9_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_nl;
  wire[6:0] FpAdd_6U_10U_7_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_7_is_a_greater_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_7_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_7_is_a_greater_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_7_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_7_is_a_greater_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_7_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_7_is_a_greater_acc_nl;
  wire[6:0] FpAdd_6U_10U_6_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_6_is_a_greater_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_6_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_6_is_a_greater_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_6_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_6_is_a_greater_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_6_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_6_is_a_greater_acc_nl;
  wire[6:0] FpAdd_6U_10U_5_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_5_is_a_greater_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_5_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_5_is_a_greater_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_5_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_5_is_a_greater_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_5_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_5_is_a_greater_acc_nl;
  wire[6:0] FpAdd_6U_10U_4_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_4_is_a_greater_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_4_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_4_is_a_greater_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_4_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_4_is_a_greater_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_4_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_4_is_a_greater_acc_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_nl;
  wire[5:0] o_col0_1_FpNormalize_6U_23U_4_else_acc_nl;
  wire[7:0] nl_o_col0_1_FpNormalize_6U_23U_4_else_acc_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[6:0] nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_4_nl;
  wire[0:0] FpAdd_6U_10U_4_and_5_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_2_nl;
  wire[5:0] o_col0_2_FpNormalize_6U_23U_4_else_acc_nl;
  wire[7:0] nl_o_col0_2_FpNormalize_6U_23U_4_else_acc_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[6:0] nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_10_nl;
  wire[0:0] FpAdd_6U_10U_4_and_11_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_4_nl;
  wire[5:0] o_col0_3_FpNormalize_6U_23U_4_else_acc_nl;
  wire[7:0] nl_o_col0_3_FpNormalize_6U_23U_4_else_acc_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[6:0] nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_16_nl;
  wire[0:0] FpAdd_6U_10U_4_and_17_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_6_nl;
  wire[5:0] o_col0_4_FpNormalize_6U_23U_4_else_acc_nl;
  wire[7:0] nl_o_col0_4_FpNormalize_6U_23U_4_else_acc_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[6:0] nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_and_22_nl;
  wire[0:0] FpAdd_6U_10U_4_and_23_nl;
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_nl;
  wire[5:0] o_col1_1_FpNormalize_6U_23U_5_else_acc_nl;
  wire[7:0] nl_o_col1_1_FpNormalize_6U_23U_5_else_acc_nl;
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[6:0] nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_4_nl;
  wire[0:0] FpAdd_6U_10U_5_and_5_nl;
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_2_nl;
  wire[5:0] o_col1_2_FpNormalize_6U_23U_5_else_acc_nl;
  wire[7:0] nl_o_col1_2_FpNormalize_6U_23U_5_else_acc_nl;
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[6:0] nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_10_nl;
  wire[0:0] FpAdd_6U_10U_5_and_11_nl;
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_4_nl;
  wire[5:0] o_col1_3_FpNormalize_6U_23U_5_else_acc_nl;
  wire[7:0] nl_o_col1_3_FpNormalize_6U_23U_5_else_acc_nl;
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[6:0] nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_16_nl;
  wire[0:0] FpAdd_6U_10U_5_and_17_nl;
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl;
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_6_nl;
  wire[5:0] o_col1_4_FpNormalize_6U_23U_5_else_acc_nl;
  wire[7:0] nl_o_col1_4_FpNormalize_6U_23U_5_else_acc_nl;
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[6:0] nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_5_and_22_nl;
  wire[0:0] FpAdd_6U_10U_5_and_23_nl;
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_nl;
  wire[5:0] o_col2_1_FpNormalize_6U_23U_6_else_acc_nl;
  wire[7:0] nl_o_col2_1_FpNormalize_6U_23U_6_else_acc_nl;
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[6:0] nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_4_nl;
  wire[0:0] FpAdd_6U_10U_6_and_5_nl;
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_2_nl;
  wire[5:0] o_col2_2_FpNormalize_6U_23U_6_else_acc_nl;
  wire[7:0] nl_o_col2_2_FpNormalize_6U_23U_6_else_acc_nl;
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[6:0] nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_10_nl;
  wire[0:0] FpAdd_6U_10U_6_and_11_nl;
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_4_nl;
  wire[5:0] o_col2_3_FpNormalize_6U_23U_6_else_acc_nl;
  wire[7:0] nl_o_col2_3_FpNormalize_6U_23U_6_else_acc_nl;
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[6:0] nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_16_nl;
  wire[0:0] FpAdd_6U_10U_6_and_17_nl;
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl;
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_6_nl;
  wire[5:0] o_col2_4_FpNormalize_6U_23U_6_else_acc_nl;
  wire[7:0] nl_o_col2_4_FpNormalize_6U_23U_6_else_acc_nl;
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[6:0] nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_6_and_22_nl;
  wire[0:0] FpAdd_6U_10U_6_and_23_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_nl;
  wire[5:0] o_col3_1_FpNormalize_6U_23U_7_else_acc_nl;
  wire[7:0] nl_o_col3_1_FpNormalize_6U_23U_7_else_acc_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[6:0] nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_4_nl;
  wire[0:0] FpAdd_6U_10U_7_and_5_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_2_nl;
  wire[5:0] o_col3_2_FpNormalize_6U_23U_7_else_acc_nl;
  wire[7:0] nl_o_col3_2_FpNormalize_6U_23U_7_else_acc_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[6:0] nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_10_nl;
  wire[0:0] FpAdd_6U_10U_7_and_11_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_4_nl;
  wire[5:0] o_col3_3_FpNormalize_6U_23U_7_else_acc_nl;
  wire[7:0] nl_o_col3_3_FpNormalize_6U_23U_7_else_acc_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[6:0] nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_16_nl;
  wire[0:0] FpAdd_6U_10U_7_and_17_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[6:0] nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[6:0] nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl;
  wire[5:0] FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_6_nl;
  wire[5:0] o_col3_4_FpNormalize_6U_23U_7_else_acc_nl;
  wire[7:0] nl_o_col3_4_FpNormalize_6U_23U_7_else_acc_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[6:0] nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_and_22_nl;
  wire[0:0] FpAdd_6U_10U_7_and_23_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_165_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_253_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_154_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_251_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_143_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_249_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_132_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_247_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_121_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_245_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_110_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_243_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_99_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_241_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_88_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_239_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_77_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_237_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_66_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_235_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_55_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_233_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_44_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_231_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_33_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_229_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_22_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_227_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_11_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_225_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl;
  wire[9:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_nl;
  wire[0:0] FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_223_nl;
  wire[0:0] data_truncate_1_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_2_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_3_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_4_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_5_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_6_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_7_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_8_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_9_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_10_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_11_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_12_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_13_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_14_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_15_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] data_truncate_16_FpMantDecShiftRight_10U_6U_10U_carry_and_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_15_nl;
  wire[0:0] FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_3_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_15_nl;
  wire[0:0] FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_3_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_15_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_3_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl;
  wire[0:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_3_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl;
  wire[9:0] m_row0_4_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_m_row0_4_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl;
  wire[9:0] m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_3_nl;
  wire[9:0] m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[10:0] nl_m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_3_nl;
  wire[9:0] m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[10:0] nl_m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_nl;
  wire[0:0] FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_1_nl;
  wire[0:0] FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_2_nl;
  wire[0:0] FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_3_nl;
  wire[0:0] FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_nl;
  wire[0:0] FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_1_nl;
  wire[0:0] FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_2_nl;
  wire[0:0] FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_3_nl;
  wire[0:0] FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_nl;
  wire[0:0] FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_1_nl;
  wire[0:0] FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_2_nl;
  wire[0:0] FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_3_nl;
  wire[0:0] FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_nl;
  wire[0:0] FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_1_nl;
  wire[0:0] FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_2_nl;
  wire[0:0] FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_3_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_or_9_nl;
  wire[0:0] FpAdd_6U_10U_o_sign_or_6_nl;
  wire[0:0] m_row1_if_d2_or_9_nl;
  wire[0:0] m_row1_if_d2_or_6_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_15_nl;
  wire[0:0] FpAdd_6U_10U_1_o_sign_or_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_nl;
  wire[6:0] m_row0_1_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_m_row0_1_FpNormalize_6U_23U_acc_nl;
  wire[6:0] m_row0_2_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_m_row0_2_FpNormalize_6U_23U_acc_nl;
  wire[6:0] m_row0_3_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_m_row0_3_FpNormalize_6U_23U_acc_nl;
  wire[6:0] m_row0_4_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_m_row0_4_FpNormalize_6U_23U_acc_nl;
  wire[6:0] m_row1_1_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_m_row1_1_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] m_row1_2_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_m_row1_2_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] m_row1_3_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_m_row1_3_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] m_row1_4_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_m_row1_4_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] m_row2_1_FpNormalize_6U_23U_2_acc_nl;
  wire[8:0] nl_m_row2_1_FpNormalize_6U_23U_2_acc_nl;
  wire[6:0] m_row2_2_FpNormalize_6U_23U_2_acc_nl;
  wire[8:0] nl_m_row2_2_FpNormalize_6U_23U_2_acc_nl;
  wire[6:0] m_row2_3_FpNormalize_6U_23U_2_acc_nl;
  wire[8:0] nl_m_row2_3_FpNormalize_6U_23U_2_acc_nl;
  wire[6:0] m_row2_4_FpNormalize_6U_23U_2_acc_nl;
  wire[8:0] nl_m_row2_4_FpNormalize_6U_23U_2_acc_nl;
  wire[6:0] m_row3_1_FpNormalize_6U_23U_3_acc_nl;
  wire[8:0] nl_m_row3_1_FpNormalize_6U_23U_3_acc_nl;
  wire[6:0] m_row3_2_FpNormalize_6U_23U_3_acc_nl;
  wire[8:0] nl_m_row3_2_FpNormalize_6U_23U_3_acc_nl;
  wire[6:0] m_row3_3_FpNormalize_6U_23U_3_acc_nl;
  wire[8:0] nl_m_row3_3_FpNormalize_6U_23U_3_acc_nl;
  wire[6:0] m_row3_4_FpNormalize_6U_23U_3_acc_nl;
  wire[8:0] nl_m_row3_4_FpNormalize_6U_23U_3_acc_nl;
  wire[6:0] o_col0_1_FpNormalize_6U_23U_4_acc_nl;
  wire[8:0] nl_o_col0_1_FpNormalize_6U_23U_4_acc_nl;
  wire[6:0] o_col0_2_FpNormalize_6U_23U_4_acc_nl;
  wire[8:0] nl_o_col0_2_FpNormalize_6U_23U_4_acc_nl;
  wire[6:0] o_col0_3_FpNormalize_6U_23U_4_acc_nl;
  wire[8:0] nl_o_col0_3_FpNormalize_6U_23U_4_acc_nl;
  wire[6:0] o_col0_4_FpNormalize_6U_23U_4_acc_nl;
  wire[8:0] nl_o_col0_4_FpNormalize_6U_23U_4_acc_nl;
  wire[6:0] o_col1_1_FpNormalize_6U_23U_5_acc_nl;
  wire[8:0] nl_o_col1_1_FpNormalize_6U_23U_5_acc_nl;
  wire[6:0] o_col1_2_FpNormalize_6U_23U_5_acc_nl;
  wire[8:0] nl_o_col1_2_FpNormalize_6U_23U_5_acc_nl;
  wire[6:0] o_col1_3_FpNormalize_6U_23U_5_acc_nl;
  wire[8:0] nl_o_col1_3_FpNormalize_6U_23U_5_acc_nl;
  wire[6:0] o_col1_4_FpNormalize_6U_23U_5_acc_nl;
  wire[8:0] nl_o_col1_4_FpNormalize_6U_23U_5_acc_nl;
  wire[6:0] o_col2_1_FpNormalize_6U_23U_6_acc_nl;
  wire[8:0] nl_o_col2_1_FpNormalize_6U_23U_6_acc_nl;
  wire[6:0] o_col2_2_FpNormalize_6U_23U_6_acc_nl;
  wire[8:0] nl_o_col2_2_FpNormalize_6U_23U_6_acc_nl;
  wire[6:0] o_col2_3_FpNormalize_6U_23U_6_acc_nl;
  wire[8:0] nl_o_col2_3_FpNormalize_6U_23U_6_acc_nl;
  wire[6:0] o_col2_4_FpNormalize_6U_23U_6_acc_nl;
  wire[8:0] nl_o_col2_4_FpNormalize_6U_23U_6_acc_nl;
  wire[6:0] o_col3_1_FpNormalize_6U_23U_7_acc_nl;
  wire[8:0] nl_o_col3_1_FpNormalize_6U_23U_7_acc_nl;
  wire[6:0] o_col3_2_FpNormalize_6U_23U_7_acc_nl;
  wire[8:0] nl_o_col3_2_FpNormalize_6U_23U_7_acc_nl;
  wire[6:0] o_col3_3_FpNormalize_6U_23U_7_acc_nl;
  wire[8:0] nl_o_col3_3_FpNormalize_6U_23U_7_acc_nl;
  wire[6:0] o_col3_4_FpNormalize_6U_23U_7_acc_nl;
  wire[8:0] nl_o_col3_4_FpNormalize_6U_23U_7_acc_nl;
  wire[0:0] or_92_nl;
  wire[0:0] or_102_nl;
  wire[0:0] or_112_nl;
  wire[0:0] or_127_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] or_145_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] or_163_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] or_176_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] or_310_nl;
  wire[0:0] or_323_nl;
  wire[0:0] or_340_nl;
  wire[0:0] or_357_nl;
  wire[0:0] or_380_nl;
  wire[0:0] or_397_nl;
  wire[0:0] or_414_nl;
  wire[0:0] or_440_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] or_454_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] or_462_nl;
  wire[0:0] or_486_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] or_500_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] or_506_nl;
  wire[0:0] and_2496_nl;
  wire[0:0] or_534_nl;
  wire[0:0] or_553_nl;
  wire[0:0] or_572_nl;
  wire[0:0] or_600_nl;
  wire[0:0] or_620_nl;
  wire[0:0] and_2636_nl;
  wire[0:0] or_626_nl;
  wire[0:0] and_2634_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] and_2457_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] and_2458_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] and_2449_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] and_2450_nl;
  wire[0:0] or_843_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] or_1226_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] mux_660_nl;
  wire[10:0] FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl;
  wire[10:0] FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl;
  wire[10:0] FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl;
  wire[10:0] FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl;
  wire[10:0] FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl;
  wire[10:0] FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl;
  wire[10:0] FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl;
  wire[10:0] FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_160_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_161_nl;
  wire[0:0] data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_162_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_163_nl;
  wire[0:0] data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_164_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_165_nl;
  wire[0:0] data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_166_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_167_nl;
  wire[0:0] data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_168_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_169_nl;
  wire[0:0] data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_170_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_171_nl;
  wire[0:0] data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_172_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_173_nl;
  wire[0:0] data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_174_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_175_nl;
  wire[0:0] data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_176_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_177_nl;
  wire[0:0] data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_178_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_179_nl;
  wire[0:0] data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_180_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_181_nl;
  wire[0:0] data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_182_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_183_nl;
  wire[0:0] data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_184_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_185_nl;
  wire[0:0] data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_186_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_187_nl;
  wire[0:0] data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_188_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_189_nl;
  wire[0:0] data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;
  wire[17:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_190_nl;
  wire[0:0] IntShiftRight_18U_2U_8U_obits_fixed_mux_191_nl;
  wire[0:0] data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl;
  wire[0:0] data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [8:0] nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a;
  assign nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[136:128];
  wire [5:0] nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s;
  assign nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_33)
      + 5'b1;
  wire [8:0] nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[8:0];
  wire [5:0] nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_32)
      + 5'b1;
  wire [8:0] nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a;
  assign nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[152:144];
  wire [5:0] nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s;
  assign nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_35)
      + 5'b1;
  wire [8:0] nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[24:16];
  wire [5:0] nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_34)
      + 5'b1;
  wire [8:0] nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a;
  assign nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[168:160];
  wire [5:0] nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s;
  assign nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_37)
      + 5'b1;
  wire [8:0] nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[40:32];
  wire [5:0] nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_36)
      + 5'b1;
  wire [10:0] nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a = {m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_is_a_greater_oelse_not_33_nl;
  wire [7:0] nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2}) + ({(~ (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]))
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = nl_m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_3_is_a_greater_oelse_not_33_nl = ~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp;
  assign m_row3_4_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_4_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_3_is_a_greater_oelse_not_33_nl)));
  assign nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_4_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row3_4_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl;
  wire [10:0] nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a;
  assign m_row3_4_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a = {(m_row3_4_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2)}) + 6'b1;
  assign m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = nl_m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl[5:0];
  assign m_row3_4_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_4_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp));
  assign nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_4_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [8:0] nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[104:96];
  wire [5:0] nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_42)
      + 5'b1;
  wire [8:0] nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a;
  assign nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[232:224];
  wire [5:0] nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s;
  assign nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_46)
      + 5'b1;
  wire [10:0] nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a = {m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_is_a_greater_oelse_not_30_nl;
  wire [7:0] nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = nl_m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_3_is_a_greater_oelse_not_30_nl = ~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp;
  assign m_row3_3_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_3_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_3_is_a_greater_oelse_not_30_nl)));
  assign nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_3_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row3_3_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl;
  wire [10:0] nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a;
  assign m_row3_3_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a = {(m_row3_3_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = nl_m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl[5:0];
  assign m_row3_3_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_3_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp));
  assign nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_3_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [8:0] nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[88:80];
  wire [5:0] nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_41)
      + 5'b1;
  wire [8:0] nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a;
  assign nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[216:208];
  wire [5:0] nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s;
  assign nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_45)
      + 5'b1;
  wire [10:0] nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a = {m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = nl_m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_3_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp;
  assign m_row3_2_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_2_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_3_is_a_greater_oelse_not_27_nl)));
  assign nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_2_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row3_2_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl;
  wire [10:0] nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a;
  assign m_row3_2_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a = {(m_row3_2_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = nl_m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl[5:0];
  assign m_row3_2_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_2_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp));
  assign nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_2_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [8:0] nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[72:64];
  wire [5:0] nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_40)
      + 5'b1;
  wire [8:0] nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a;
  assign nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[200:192];
  wire [5:0] nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s;
  assign nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_44)
      + 5'b1;
  wire [10:0] nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a = {m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_3_is_a_greater_oelse_not_24_nl;
  wire [7:0] nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl = nl_m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_3_is_a_greater_oelse_not_24_nl = ~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp;
  assign m_row3_1_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_1_FpAdd_6U_10U_3_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_3_is_a_greater_oelse_not_24_nl)));
  assign nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_1_FpAdd_6U_10U_3_a_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row3_1_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl;
  wire [10:0] nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a;
  assign m_row3_1_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a = {(m_row3_1_FpAdd_6U_10U_3_IsZero_6U_10U_7_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0};
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl;
  wire[5:0] m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl = nl_m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl[5:0];
  assign m_row3_1_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row3_1_FpAdd_6U_10U_3_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp));
  assign nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row3_1_FpAdd_6U_10U_3_b_left_shift_FpAdd_6U_10U_3_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a = {m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1};
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_is_a_greater_oelse_not_33_nl;
  wire [7:0] nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]))
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = nl_m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_2_is_a_greater_oelse_not_33_nl = ~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp;
  assign m_row2_4_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_4_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_2_is_a_greater_oelse_not_33_nl)));
  assign nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_4_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a = {m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0};
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]))
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = nl_m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl[5:0];
  assign m_row2_4_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_4_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp));
  assign nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_4_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a = {m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_7_cse};
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_is_a_greater_oelse_not_30_nl;
  wire [7:0] nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = nl_m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_2_is_a_greater_oelse_not_30_nl = ~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp;
  assign m_row2_3_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_3_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_2_is_a_greater_oelse_not_30_nl)));
  assign nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_3_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a = {m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0};
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = nl_m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl[5:0];
  assign m_row2_3_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_3_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp));
  assign nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_3_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a = {m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_4_cse};
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = nl_m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_2_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp;
  assign m_row2_2_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_2_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_2_is_a_greater_oelse_not_27_nl)));
  assign nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_2_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a = {m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0};
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = nl_m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl[5:0];
  assign m_row2_2_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_2_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp));
  assign nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_2_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a = {m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_1_cse};
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_2_is_a_greater_oelse_not_24_nl;
  wire [7:0] nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl = nl_m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_2_is_a_greater_oelse_not_24_nl = ~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp;
  assign m_row2_1_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_1_FpAdd_6U_10U_2_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_2_is_a_greater_oelse_not_24_nl)));
  assign nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_1_FpAdd_6U_10U_2_a_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a = {m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0};
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl;
  wire[5:0] m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl = nl_m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl[5:0];
  assign m_row2_1_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row2_1_FpAdd_6U_10U_2_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp));
  assign nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row2_1_FpAdd_6U_10U_2_b_left_shift_FpAdd_6U_10U_2_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row1_4_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl;
  wire [10:0] nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign m_row1_4_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl = ~(m_row2_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {(m_row1_4_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0};
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_33_nl;
  wire [7:0] nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_33_nl = ~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp;
  assign m_row1_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_33_nl)));
  assign nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1};
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]))
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign m_row1_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp));
  assign nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row1_3_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl;
  wire [10:0] nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign m_row1_3_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl = ~(m_row2_3_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {(m_row1_3_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0};
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_30_nl;
  wire [7:0] nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)})
      + 6'b1;
  assign m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_30_nl = ~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp;
  assign m_row1_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_30_nl)));
  assign nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_7_cse};
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign m_row1_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp));
  assign nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row1_2_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl;
  wire [10:0] nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign m_row1_2_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl = ~(m_row2_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {(m_row1_2_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0};
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)})
      + 6'b1;
  assign m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp;
  assign m_row1_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl)));
  assign nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_4_cse};
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign m_row1_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp));
  assign nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row1_1_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl;
  wire [10:0] nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign m_row1_1_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl = ~(m_row2_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {(m_row1_1_FpAdd_6U_10U_1_IsZero_6U_10U_2_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0};
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_24_nl;
  wire [7:0] nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)})
      + 6'b1;
  assign m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_24_nl = ~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp;
  assign m_row1_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_24_nl)));
  assign nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10
      , m_row2_if_d1_mux_1_cse};
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign m_row1_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (m_row1_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp));
  assign nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row1_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_nand_nl;
  wire [10:0] nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {(m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0};
  wire[5:0] m_row0_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_33_nl;
  wire [7:0] nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2)}) + 6'b1;
  assign m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = nl_m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_is_a_greater_oelse_not_33_nl = ~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp;
  assign m_row0_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_4_FpAdd_6U_10U_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_is_a_greater_oelse_not_33_nl)));
  assign nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl;
  wire [10:0] nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl = ~(m_row1_4_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {(m_row0_4_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1};
  wire[5:0] m_row0_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl = nl_m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl[5:0];
  assign m_row0_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_4_FpAdd_6U_10U_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp));
  assign nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_nand_nl;
  wire [10:0] nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {(m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0};
  wire[5:0] m_row0_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_30_nl;
  wire [7:0] nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = nl_m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_is_a_greater_oelse_not_30_nl = ~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp;
  assign m_row0_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_3_FpAdd_6U_10U_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_is_a_greater_oelse_not_30_nl)));
  assign nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl;
  wire [10:0] nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl = ~(m_row1_3_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {(m_row0_3_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl)
      , m_row2_if_d1_mux_7_cse};
  wire[5:0] m_row0_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl = nl_m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl[5:0];
  assign m_row0_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_3_FpAdd_6U_10U_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp));
  assign nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_nand_nl;
  wire [10:0] nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {(m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0};
  wire[5:0] m_row0_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = nl_m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp;
  assign m_row0_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_2_FpAdd_6U_10U_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_is_a_greater_oelse_not_27_nl)));
  assign nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl;
  wire [10:0] nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl = ~(m_row1_2_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {(m_row0_2_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl)
      , m_row2_if_d1_mux_4_cse};
  wire[5:0] m_row0_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl = nl_m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl[5:0];
  assign m_row0_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_2_FpAdd_6U_10U_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp));
  assign nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_nand_nl;
  wire [10:0] nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_nand_nl = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0==10'b0000000000)
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2!=4'b0000))));
  assign nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {(m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_nand_nl)
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0};
  wire[5:0] m_row0_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_24_nl;
  wire [7:0] nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + ({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2)})
      + 6'b1;
  assign m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl = nl_m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_is_a_greater_oelse_not_24_nl = ~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp;
  assign m_row0_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_1_FpAdd_6U_10U_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_is_a_greater_oelse_not_24_nl)));
  assign nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire[0:0] m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl;
  wire [10:0] nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl = ~(m_row1_1_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4!=2'b00) | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {(m_row0_1_FpAdd_6U_10U_IsZero_6U_10U_1_nand_nl)
      , m_row2_if_d1_mux_1_cse};
  wire[5:0] m_row0_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire[7:0] nl_m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl;
  wire [7:0] nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign nl_m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3
      , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2}) + ({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 6'b1;
  assign m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl = nl_m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl[5:0];
  assign m_row0_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl =
      ~(MUX_v_6_2_2(6'b000000, (m_row0_1_FpAdd_6U_10U_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp));
  assign nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (m_row0_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [8:0] nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a;
  assign nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[184:176];
  wire [5:0] nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s;
  assign nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_39)
      + 5'b1;
  wire [8:0] nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[56:48];
  wire [5:0] nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_38)
      + 5'b1;
  wire [8:0] nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[120:112];
  wire [5:0] nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_43)
      + 5'b1;
  wire [8:0] nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a;
  assign nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a = chn_data_in_rsci_d_mxwt[248:240];
  wire [5:0] nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s;
  assign nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_47)
      + 5'b1;
  wire[17:0] o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire[18:0] nl_o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire [20:0] nl_data_truncate_16_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_2_o_acc_2_itm_2)
      + conv_s2s_17_18(m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2);
  assign o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl = nl_o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl[17:0];
  assign nl_data_truncate_16_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col3_4_IntSubExt_17U_17U_18U_2_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire[18:0] nl_o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire [20:0] nl_data_truncate_15_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl = conv_s2s_17_18(m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2)
      - conv_s2s_17_18(m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2);
  assign o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl = nl_o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl[17:0];
  assign nl_data_truncate_15_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col2_4_IntSubExt_17U_17U_18U_1_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl;
  wire[18:0] nl_o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl;
  wire [20:0] nl_data_truncate_14_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl = conv_s2s_17_18(m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2)
      + conv_s2s_17_18(m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2);
  assign o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl = nl_o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl[17:0];
  assign nl_data_truncate_14_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col1_4_IntAddExt_17U_17U_18U_o_acc_nl)
      , 3'b0};
  wire[17:0] IntSubExt_16U_16U_17U_2_o_acc_nl;
  wire[18:0] nl_IntSubExt_16U_16U_17U_2_o_acc_nl;
  wire [20:0] nl_data_truncate_13_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_IntSubExt_16U_16U_17U_2_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_2_o_acc_1_itm_2)
      - conv_s2s_17_18(m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2);
  assign IntSubExt_16U_16U_17U_2_o_acc_nl = nl_IntSubExt_16U_16U_17U_2_o_acc_nl[17:0];
  assign nl_data_truncate_13_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(IntSubExt_16U_16U_17U_2_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire[18:0] nl_o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire [20:0] nl_data_truncate_12_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_1_o_acc_2_itm_2)
      + conv_s2s_17_18(m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2);
  assign o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl = nl_o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl[17:0];
  assign nl_data_truncate_12_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col3_3_IntSubExt_17U_17U_18U_2_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire[18:0] nl_o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire [20:0] nl_data_truncate_11_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl = conv_s2s_17_18(m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2)
      - conv_s2s_17_18(m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2);
  assign o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl = nl_o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl[17:0];
  assign nl_data_truncate_11_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col2_3_IntSubExt_17U_17U_18U_1_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl;
  wire[18:0] nl_o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl;
  wire [20:0] nl_data_truncate_10_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl = conv_s2s_17_18(m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2)
      + conv_s2s_17_18(m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2);
  assign o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl = nl_o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl[17:0];
  assign nl_data_truncate_10_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col1_3_IntAddExt_17U_17U_18U_o_acc_nl)
      , 3'b0};
  wire[17:0] IntSubExt_16U_16U_17U_1_o_acc_nl;
  wire[18:0] nl_IntSubExt_16U_16U_17U_1_o_acc_nl;
  wire [20:0] nl_data_truncate_9_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_IntSubExt_16U_16U_17U_1_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_1_o_acc_1_itm_2)
      - conv_s2s_17_18(m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2);
  assign IntSubExt_16U_16U_17U_1_o_acc_nl = nl_IntSubExt_16U_16U_17U_1_o_acc_nl[17:0];
  assign nl_data_truncate_9_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(IntSubExt_16U_16U_17U_1_o_acc_nl)
      , 3'b0};
  wire[17:0] IntAddExt_16U_16U_17U_o_acc_2_nl;
  wire[19:0] nl_IntAddExt_16U_16U_17U_o_acc_2_nl;
  wire [20:0] nl_data_truncate_8_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_IntAddExt_16U_16U_17U_o_acc_2_nl = conv_s2s_17_18(IntAddExt_16U_16U_17U_o_acc_1_itm_2)
      + conv_s2s_17_18(m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2) + 18'b1;
  assign IntAddExt_16U_16U_17U_o_acc_2_nl = nl_IntAddExt_16U_16U_17U_o_acc_2_nl[17:0];
  assign nl_data_truncate_8_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(IntAddExt_16U_16U_17U_o_acc_2_nl)
      , 3'b0};
  wire[17:0] o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire[18:0] nl_o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire [20:0] nl_data_truncate_7_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl = conv_s2s_17_18(m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2)
      - conv_s2s_17_18(m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl = nl_o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl[17:0];
  assign nl_data_truncate_7_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col2_2_IntSubExt_17U_17U_18U_1_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl;
  wire[18:0] nl_o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl;
  wire [20:0] nl_data_truncate_6_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl = conv_s2s_17_18(m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2)
      + conv_s2s_17_18(m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl = nl_o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl[17:0];
  assign nl_data_truncate_6_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col1_2_IntAddExt_17U_17U_18U_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl;
  wire[18:0] nl_o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl;
  wire [20:0] nl_data_truncate_5_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl = conv_s2s_17_18(IntAddExt_16U_16U_17U_o_acc_itm_2)
      + conv_s2s_17_18(~ m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl = nl_o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl[17:0];
  assign nl_data_truncate_5_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col0_2_IntSubExt_17U_17U_18U_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire[18:0] nl_o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl;
  wire [20:0] nl_data_truncate_4_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_o_acc_2_itm_2)
      + conv_s2s_17_18(m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl = nl_o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl[17:0];
  assign nl_data_truncate_4_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col3_1_IntSubExt_17U_17U_18U_2_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire[18:0] nl_o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl;
  wire [20:0] nl_data_truncate_3_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl = conv_s2s_17_18(m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2)
      - conv_s2s_17_18(m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl = nl_o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl[17:0];
  assign nl_data_truncate_3_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col2_1_IntSubExt_17U_17U_18U_1_o_acc_nl)
      , 3'b0};
  wire[17:0] o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl;
  wire[18:0] nl_o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl;
  wire [20:0] nl_data_truncate_2_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl = conv_s2s_17_18(m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2)
      + conv_s2s_17_18(m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl = nl_o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl[17:0];
  assign nl_data_truncate_2_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(o_col1_1_IntAddExt_17U_17U_18U_o_acc_nl)
      , 3'b0};
  wire[17:0] IntSubExt_16U_16U_17U_o_acc_nl;
  wire[18:0] nl_IntSubExt_16U_16U_17U_o_acc_nl;
  wire [20:0] nl_data_truncate_1_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a;
  assign nl_IntSubExt_16U_16U_17U_o_acc_nl = conv_s2s_17_18(IntSubExt_16U_16U_17U_o_acc_1_itm_2)
      - conv_s2s_17_18(m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2);
  assign IntSubExt_16U_16U_17U_o_acc_nl = nl_IntSubExt_16U_16U_17U_o_acc_nl[17:0];
  assign nl_data_truncate_1_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a = {(IntSubExt_16U_16U_17U_o_acc_nl)
      , 3'b0};
  wire [9:0] nl_m_row0_1_leading_sign_10_0_rg_mantissa;
  assign nl_m_row0_1_leading_sign_10_0_rg_mantissa = chn_data_in_rsci_d_mxwt[9:0];
  wire [9:0] nl_m_row0_1_leading_sign_10_0_1_rg_mantissa;
  assign nl_m_row0_1_leading_sign_10_0_1_rg_mantissa = chn_data_in_rsci_d_mxwt[137:128];
  wire [9:0] nl_m_row0_2_leading_sign_10_0_rg_mantissa;
  assign nl_m_row0_2_leading_sign_10_0_rg_mantissa = chn_data_in_rsci_d_mxwt[25:16];
  wire [9:0] nl_m_row0_2_leading_sign_10_0_1_rg_mantissa;
  assign nl_m_row0_2_leading_sign_10_0_1_rg_mantissa = chn_data_in_rsci_d_mxwt[153:144];
  wire [9:0] nl_m_row0_3_leading_sign_10_0_rg_mantissa;
  assign nl_m_row0_3_leading_sign_10_0_rg_mantissa = chn_data_in_rsci_d_mxwt[41:32];
  wire [9:0] nl_m_row0_3_leading_sign_10_0_1_rg_mantissa;
  assign nl_m_row0_3_leading_sign_10_0_1_rg_mantissa = chn_data_in_rsci_d_mxwt[169:160];
  wire [9:0] nl_m_row0_4_leading_sign_10_0_rg_mantissa;
  assign nl_m_row0_4_leading_sign_10_0_rg_mantissa = chn_data_in_rsci_d_mxwt[57:48];
  wire [9:0] nl_m_row0_4_leading_sign_10_0_1_rg_mantissa;
  assign nl_m_row0_4_leading_sign_10_0_1_rg_mantissa = chn_data_in_rsci_d_mxwt[185:176];
  wire [9:0] nl_m_row1_1_leading_sign_10_0_2_rg_mantissa;
  assign nl_m_row1_1_leading_sign_10_0_2_rg_mantissa = chn_data_in_rsci_d_mxwt[73:64];
  wire [9:0] nl_m_row1_2_leading_sign_10_0_2_rg_mantissa;
  assign nl_m_row1_2_leading_sign_10_0_2_rg_mantissa = chn_data_in_rsci_d_mxwt[89:80];
  wire [9:0] nl_m_row1_3_leading_sign_10_0_2_rg_mantissa;
  assign nl_m_row1_3_leading_sign_10_0_2_rg_mantissa = chn_data_in_rsci_d_mxwt[105:96];
  wire [9:0] nl_m_row1_4_leading_sign_10_0_2_rg_mantissa;
  assign nl_m_row1_4_leading_sign_10_0_2_rg_mantissa = chn_data_in_rsci_d_mxwt[121:112];
  wire [9:0] nl_m_row3_1_leading_sign_10_0_7_rg_mantissa;
  assign nl_m_row3_1_leading_sign_10_0_7_rg_mantissa = chn_data_in_rsci_d_mxwt[201:192];
  wire [9:0] nl_m_row3_2_leading_sign_10_0_7_rg_mantissa;
  assign nl_m_row3_2_leading_sign_10_0_7_rg_mantissa = chn_data_in_rsci_d_mxwt[217:208];
  wire [9:0] nl_m_row3_3_leading_sign_10_0_7_rg_mantissa;
  assign nl_m_row3_3_leading_sign_10_0_7_rg_mantissa = chn_data_in_rsci_d_mxwt[233:224];
  wire [9:0] nl_m_row3_4_leading_sign_10_0_7_rg_mantissa;
  assign nl_m_row3_4_leading_sign_10_0_7_rg_mantissa = chn_data_in_rsci_d_mxwt[249:240];
  wire [22:0] nl_o_col0_1_FpNormalize_6U_23U_4_else_lshift_rg_a;
  assign nl_o_col0_1_FpNormalize_6U_23U_4_else_lshift_rg_a = FpAdd_6U_10U_4_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col0_1_leading_sign_23_0_4_rg_mantissa;
  assign nl_o_col0_1_leading_sign_23_0_4_rg_mantissa = FpAdd_6U_10U_4_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col0_2_FpNormalize_6U_23U_4_else_lshift_rg_a;
  assign nl_o_col0_2_FpNormalize_6U_23U_4_else_lshift_rg_a = FpAdd_6U_10U_4_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col0_2_leading_sign_23_0_4_rg_mantissa;
  assign nl_o_col0_2_leading_sign_23_0_4_rg_mantissa = FpAdd_6U_10U_4_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col0_3_FpNormalize_6U_23U_4_else_lshift_rg_a;
  assign nl_o_col0_3_FpNormalize_6U_23U_4_else_lshift_rg_a = FpAdd_6U_10U_4_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col0_3_leading_sign_23_0_4_rg_mantissa;
  assign nl_o_col0_3_leading_sign_23_0_4_rg_mantissa = FpAdd_6U_10U_4_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col0_4_FpNormalize_6U_23U_4_else_lshift_rg_a;
  assign nl_o_col0_4_FpNormalize_6U_23U_4_else_lshift_rg_a = FpAdd_6U_10U_4_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col0_4_leading_sign_23_0_4_rg_mantissa;
  assign nl_o_col0_4_leading_sign_23_0_4_rg_mantissa = FpAdd_6U_10U_4_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col1_1_FpNormalize_6U_23U_5_else_lshift_rg_a;
  assign nl_o_col1_1_FpNormalize_6U_23U_5_else_lshift_rg_a = FpAdd_6U_10U_5_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col1_1_leading_sign_23_0_5_rg_mantissa;
  assign nl_o_col1_1_leading_sign_23_0_5_rg_mantissa = FpAdd_6U_10U_5_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col1_2_FpNormalize_6U_23U_5_else_lshift_rg_a;
  assign nl_o_col1_2_FpNormalize_6U_23U_5_else_lshift_rg_a = FpAdd_6U_10U_5_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col1_2_leading_sign_23_0_5_rg_mantissa;
  assign nl_o_col1_2_leading_sign_23_0_5_rg_mantissa = FpAdd_6U_10U_5_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col1_3_FpNormalize_6U_23U_5_else_lshift_rg_a;
  assign nl_o_col1_3_FpNormalize_6U_23U_5_else_lshift_rg_a = FpAdd_6U_10U_5_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col1_3_leading_sign_23_0_5_rg_mantissa;
  assign nl_o_col1_3_leading_sign_23_0_5_rg_mantissa = FpAdd_6U_10U_5_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col1_4_FpNormalize_6U_23U_5_else_lshift_rg_a;
  assign nl_o_col1_4_FpNormalize_6U_23U_5_else_lshift_rg_a = FpAdd_6U_10U_5_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col1_4_leading_sign_23_0_5_rg_mantissa;
  assign nl_o_col1_4_leading_sign_23_0_5_rg_mantissa = FpAdd_6U_10U_5_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col2_1_FpNormalize_6U_23U_6_else_lshift_rg_a;
  assign nl_o_col2_1_FpNormalize_6U_23U_6_else_lshift_rg_a = FpAdd_6U_10U_6_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col2_1_leading_sign_23_0_6_rg_mantissa;
  assign nl_o_col2_1_leading_sign_23_0_6_rg_mantissa = FpAdd_6U_10U_6_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col2_2_FpNormalize_6U_23U_6_else_lshift_rg_a;
  assign nl_o_col2_2_FpNormalize_6U_23U_6_else_lshift_rg_a = FpAdd_6U_10U_6_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col2_2_leading_sign_23_0_6_rg_mantissa;
  assign nl_o_col2_2_leading_sign_23_0_6_rg_mantissa = FpAdd_6U_10U_6_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col2_3_FpNormalize_6U_23U_6_else_lshift_rg_a;
  assign nl_o_col2_3_FpNormalize_6U_23U_6_else_lshift_rg_a = FpAdd_6U_10U_6_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col2_3_leading_sign_23_0_6_rg_mantissa;
  assign nl_o_col2_3_leading_sign_23_0_6_rg_mantissa = FpAdd_6U_10U_6_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col2_4_FpNormalize_6U_23U_6_else_lshift_rg_a;
  assign nl_o_col2_4_FpNormalize_6U_23U_6_else_lshift_rg_a = FpAdd_6U_10U_6_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col2_4_leading_sign_23_0_6_rg_mantissa;
  assign nl_o_col2_4_leading_sign_23_0_6_rg_mantissa = FpAdd_6U_10U_6_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col3_1_FpNormalize_6U_23U_7_else_lshift_rg_a;
  assign nl_o_col3_1_FpNormalize_6U_23U_7_else_lshift_rg_a = FpAdd_6U_10U_7_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col3_1_leading_sign_23_0_7_rg_mantissa;
  assign nl_o_col3_1_leading_sign_23_0_7_rg_mantissa = FpAdd_6U_10U_7_int_mant_p1_1_sva_3[22:0];
  wire [22:0] nl_o_col3_2_FpNormalize_6U_23U_7_else_lshift_rg_a;
  assign nl_o_col3_2_FpNormalize_6U_23U_7_else_lshift_rg_a = FpAdd_6U_10U_7_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col3_2_leading_sign_23_0_7_rg_mantissa;
  assign nl_o_col3_2_leading_sign_23_0_7_rg_mantissa = FpAdd_6U_10U_7_int_mant_p1_2_sva_3[22:0];
  wire [22:0] nl_o_col3_3_FpNormalize_6U_23U_7_else_lshift_rg_a;
  assign nl_o_col3_3_FpNormalize_6U_23U_7_else_lshift_rg_a = FpAdd_6U_10U_7_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col3_3_leading_sign_23_0_7_rg_mantissa;
  assign nl_o_col3_3_leading_sign_23_0_7_rg_mantissa = FpAdd_6U_10U_7_int_mant_p1_3_sva_3[22:0];
  wire [22:0] nl_o_col3_4_FpNormalize_6U_23U_7_else_lshift_rg_a;
  assign nl_o_col3_4_FpNormalize_6U_23U_7_else_lshift_rg_a = FpAdd_6U_10U_7_int_mant_p1_sva_3[22:0];
  wire [22:0] nl_o_col3_4_leading_sign_23_0_7_rg_mantissa;
  assign nl_o_col3_4_leading_sign_23_0_7_rg_mantissa = FpAdd_6U_10U_7_int_mant_p1_sva_3[22:0];
  wire [10:0] nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_4_o_mant_1_lpi_2};
  wire [3:0] nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva , (~
      (FpAdd_6U_10U_4_o_expo_1_lpi_2[0]))};
  wire [5:0] nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva
      , (~ (FpAdd_6U_10U_4_o_expo_1_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva , (~
      (FpAdd_6U_10U_4_o_expo_1_lpi_2[0]))};
  wire [10:0] nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_5_o_mant_1_lpi_2};
  wire [3:0] nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva , (~
      (FpAdd_6U_10U_5_o_expo_1_lpi_2[0]))};
  wire [5:0] nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva
      , (~ (FpAdd_6U_10U_5_o_expo_1_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva , (~
      (FpAdd_6U_10U_5_o_expo_1_lpi_2[0]))};
  wire [10:0] nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_6_o_mant_1_lpi_2};
  wire [3:0] nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva , (~
      (FpAdd_6U_10U_6_o_expo_1_lpi_2[0]))};
  wire [5:0] nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva
      , (~ (FpAdd_6U_10U_6_o_expo_1_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva , (~
      (FpAdd_6U_10U_6_o_expo_1_lpi_2[0]))};
  wire [10:0] nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_7_o_mant_1_lpi_2};
  wire [3:0] nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva , (~
      (FpAdd_6U_10U_7_o_expo_1_lpi_2[0]))};
  wire [5:0] nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva
      , (~ (FpAdd_6U_10U_7_o_expo_1_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva , (~
      (FpAdd_6U_10U_7_o_expo_1_lpi_2[0]))};
  wire [10:0] nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_4_o_mant_2_lpi_2};
  wire [3:0] nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva , (~
      (FpAdd_6U_10U_4_o_expo_2_lpi_2[0]))};
  wire [5:0] nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva
      , (~ (FpAdd_6U_10U_4_o_expo_2_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva , (~
      (FpAdd_6U_10U_4_o_expo_2_lpi_2[0]))};
  wire [10:0] nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_5_o_mant_2_lpi_2};
  wire [3:0] nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva , (~
      (FpAdd_6U_10U_5_o_expo_2_lpi_2[0]))};
  wire [5:0] nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva
      , (~ (FpAdd_6U_10U_5_o_expo_2_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva , (~
      (FpAdd_6U_10U_5_o_expo_2_lpi_2[0]))};
  wire [10:0] nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_6_o_mant_2_lpi_2};
  wire [3:0] nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva , (~
      (FpAdd_6U_10U_6_o_expo_2_lpi_2[0]))};
  wire [5:0] nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva
      , (~ (FpAdd_6U_10U_6_o_expo_2_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva , (~
      (FpAdd_6U_10U_6_o_expo_2_lpi_2[0]))};
  wire [10:0] nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_7_o_mant_2_lpi_2};
  wire [3:0] nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva , (~
      (FpAdd_6U_10U_7_o_expo_2_lpi_2[0]))};
  wire [5:0] nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva
      , (~ (FpAdd_6U_10U_7_o_expo_2_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva , (~
      (FpAdd_6U_10U_7_o_expo_2_lpi_2[0]))};
  wire [10:0] nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a =
      {1'b1 , FpAdd_6U_10U_4_o_mant_3_lpi_2};
  wire [3:0] nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s =
      {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva , (~
      (FpAdd_6U_10U_4_o_expo_3_lpi_2[0]))};
  wire [5:0] nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva
      , (~ (FpAdd_6U_10U_4_o_expo_3_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva ,
      (~ (FpAdd_6U_10U_4_o_expo_3_lpi_2[0]))};
  wire [10:0] nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_5_o_mant_3_lpi_2};
  wire [3:0] nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva ,
      (~ (FpAdd_6U_10U_5_o_expo_3_lpi_2[0]))};
  wire [5:0] nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva
      , (~ (FpAdd_6U_10U_5_o_expo_3_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva ,
      (~ (FpAdd_6U_10U_5_o_expo_3_lpi_2[0]))};
  wire [10:0] nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_6_o_mant_3_lpi_2};
  wire [3:0] nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva ,
      (~ (FpAdd_6U_10U_6_o_expo_3_lpi_2[0]))};
  wire [5:0] nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva
      , (~ (FpAdd_6U_10U_6_o_expo_3_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva ,
      (~ (FpAdd_6U_10U_6_o_expo_3_lpi_2[0]))};
  wire [10:0] nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_7_o_mant_3_lpi_2};
  wire [3:0] nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva ,
      (~ (FpAdd_6U_10U_7_o_expo_3_lpi_2[0]))};
  wire [5:0] nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva
      , (~ (FpAdd_6U_10U_7_o_expo_3_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva ,
      (~ (FpAdd_6U_10U_7_o_expo_3_lpi_2[0]))};
  wire [10:0] nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_4_o_mant_lpi_2};
  wire [3:0] nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva ,
      (~ (FpAdd_6U_10U_4_o_expo_lpi_2[0]))};
  wire [5:0] nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva
      , (~ (FpAdd_6U_10U_4_o_expo_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva ,
      (~ (FpAdd_6U_10U_4_o_expo_lpi_2[0]))};
  wire [10:0] nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_5_o_mant_lpi_2};
  wire [3:0] nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva ,
      (~ (FpAdd_6U_10U_5_o_expo_lpi_2[0]))};
  wire [5:0] nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva
      , (~ (FpAdd_6U_10U_5_o_expo_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva ,
      (~ (FpAdd_6U_10U_5_o_expo_lpi_2[0]))};
  wire [10:0] nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_6_o_mant_lpi_2};
  wire [3:0] nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva ,
      (~ (FpAdd_6U_10U_6_o_expo_lpi_2[0]))};
  wire [5:0] nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva
      , (~ (FpAdd_6U_10U_6_o_expo_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva ,
      (~ (FpAdd_6U_10U_6_o_expo_lpi_2[0]))};
  wire [10:0] nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a;
  assign nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a
      = {1'b1 , FpAdd_6U_10U_7_o_mant_lpi_2};
  wire [3:0] nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s;
  assign nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva , (~
      (FpAdd_6U_10U_7_o_expo_lpi_2[0]))};
  wire [5:0] nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s;
  assign nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s
      = conv_u2s_4_5({FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva
      , (~ (FpAdd_6U_10U_7_o_expo_lpi_2[0]))}) + 5'b11111;
  wire [3:0] nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s;
  assign nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s
      = {FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva , (~
      (FpAdd_6U_10U_7_o_expo_lpi_2[0]))};
  wire [10:0] nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a = {reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = nl_o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl[5:0];
  assign o_col0_1_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_1_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1));
  assign nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_1_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a = {o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2
      , FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6};
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = nl_o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_4_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1;
  assign o_col0_1_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_1_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_4_is_a_greater_oelse_not_23_nl)));
  assign nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_1_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a = {reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = nl_o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl[5:0];
  assign o_col0_2_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_2_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1));
  assign nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_2_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a = {o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2
      , FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6};
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = nl_o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_4_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1;
  assign o_col0_2_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_2_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_4_is_a_greater_oelse_not_25_nl)));
  assign nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_2_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a = {reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = nl_o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl[5:0];
  assign o_col0_3_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_3_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1));
  assign nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_3_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a = {o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2
      , FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6};
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = nl_o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_4_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1;
  assign o_col0_3_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_3_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_4_is_a_greater_oelse_not_27_nl)));
  assign nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_3_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a = {reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl = nl_o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl[5:0];
  assign o_col0_4_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_4_FpAdd_6U_10U_4_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1));
  assign nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_4_FpAdd_6U_10U_4_b_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a = {o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2
      , FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6};
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl;
  wire[5:0] o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_4_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl = nl_o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_4_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1;
  assign o_col0_4_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col0_4_FpAdd_6U_10U_4_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_4_is_a_greater_oelse_not_29_nl)));
  assign nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col0_4_FpAdd_6U_10U_4_a_left_shift_FpAdd_6U_10U_4_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a = {reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire [7:0] nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s;
  assign o_col1_1_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_1_sva, FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1));
  assign nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_1_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a = {reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col1_1_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_5_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_5_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1;
  assign o_col1_1_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1, (FpAdd_6U_10U_5_is_a_greater_oelse_not_23_nl)));
  assign nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_1_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a = {reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire [7:0] nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s;
  assign o_col1_2_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_2_sva, FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1));
  assign nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_2_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a = {reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col1_2_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_5_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_5_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1;
  assign o_col1_2_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1, (FpAdd_6U_10U_5_is_a_greater_oelse_not_25_nl)));
  assign nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_2_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a = {reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire [7:0] nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s;
  assign o_col1_3_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_3_sva, FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1));
  assign nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_3_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a = {reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col1_3_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_5_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_5_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1;
  assign o_col1_3_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1, (FpAdd_6U_10U_5_is_a_greater_oelse_not_27_nl)));
  assign nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_3_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a = {reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire [7:0] nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s;
  assign o_col1_4_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_sva, FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1));
  assign nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_4_FpAdd_6U_10U_5_b_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a = {reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col1_4_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_5_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_5_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1;
  assign o_col1_4_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_sva_1, (FpAdd_6U_10U_5_is_a_greater_oelse_not_29_nl)));
  assign nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col1_4_FpAdd_6U_10U_5_a_left_shift_FpAdd_6U_10U_5_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a = {reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire [7:0] nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s;
  assign o_col2_1_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1, FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1));
  assign nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_1_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a = {reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col2_1_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_6_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_6_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1;
  assign o_col2_1_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_1_sva, (FpAdd_6U_10U_6_is_a_greater_oelse_not_23_nl)));
  assign nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_1_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a = {reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire [7:0] nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s;
  assign o_col2_2_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1, FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1));
  assign nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_2_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a = {reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1
      , FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col2_2_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_6_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_6_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1;
  assign o_col2_2_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_2_sva, (FpAdd_6U_10U_6_is_a_greater_oelse_not_25_nl)));
  assign nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_2_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a = {reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire [7:0] nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s;
  assign o_col2_3_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1, FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1));
  assign nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_3_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a = {reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col2_3_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_6_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_6_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1;
  assign o_col2_3_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_3_sva, (FpAdd_6U_10U_6_is_a_greater_oelse_not_27_nl)));
  assign nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_3_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a = {reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire [7:0] nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s;
  assign o_col2_4_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_a_right_shift_qr_sva_1, FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1));
  assign nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_4_FpAdd_6U_10U_6_b_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a = {reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse
      , FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6};
  wire[5:0] o_col2_4_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_6_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_6_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1;
  assign o_col2_4_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, FpAdd_6U_10U_5_b_right_shift_qr_sva, (FpAdd_6U_10U_6_is_a_greater_oelse_not_29_nl)));
  assign nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col2_4_FpAdd_6U_10U_6_a_left_shift_FpAdd_6U_10U_6_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a = {o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2
      , FpAdd_6U_10U_o_mant_lpi_1_dfm_6};
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = nl_o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl[5:0];
  assign o_col3_1_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_1_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1));
  assign nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_1_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a = {reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = nl_o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_7_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1;
  assign o_col3_1_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_1_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_7_is_a_greater_oelse_not_23_nl)));
  assign nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_1_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a = {o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2
      , FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6};
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = nl_o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl[5:0];
  assign o_col3_2_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_2_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1));
  assign nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_2_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a = {reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = nl_o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_7_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1;
  assign o_col3_2_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_2_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_7_is_a_greater_oelse_not_25_nl)));
  assign nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_2_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a = {o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2
      , FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6};
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = nl_o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl[5:0];
  assign o_col3_3_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_3_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1));
  assign nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_3_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a = {reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = nl_o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_7_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1;
  assign o_col3_3_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_3_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_7_is_a_greater_oelse_not_27_nl)));
  assign nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_3_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a = {o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2
      , FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6};
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire[7:0] nl_o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl;
  wire [7:0] nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl = nl_o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl[5:0];
  assign o_col3_4_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_4_FpAdd_6U_10U_7_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1));
  assign nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_4_FpAdd_6U_10U_7_b_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a;
  assign nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a = {reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse
      , FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6};
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl;
  wire[5:0] o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_7_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s;
  assign nl_o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = ({reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl = nl_o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_7_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1;
  assign o_col3_4_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (o_col3_4_FpAdd_6U_10U_7_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_7_is_a_greater_oelse_not_29_nl)));
  assign nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s = ({1'b1 , (o_col3_4_FpAdd_6U_10U_7_a_left_shift_FpAdd_6U_10U_7_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [255:0] nl_NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_inst_chn_data_out_rsci_d;
  assign nl_NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_inst_chn_data_out_rsci_d
      = {chn_data_out_rsci_d_255 , chn_data_out_rsci_d_254 , chn_data_out_rsci_d_253_250
      , chn_data_out_rsci_d_249_247 , chn_data_out_rsci_d_246_241 , chn_data_out_rsci_d_240
      , chn_data_out_rsci_d_239 , chn_data_out_rsci_d_238 , chn_data_out_rsci_d_237_234
      , chn_data_out_rsci_d_233_231 , chn_data_out_rsci_d_230_225 , chn_data_out_rsci_d_224
      , chn_data_out_rsci_d_223 , chn_data_out_rsci_d_222 , chn_data_out_rsci_d_221_218
      , chn_data_out_rsci_d_217_215 , chn_data_out_rsci_d_214_209 , chn_data_out_rsci_d_208
      , chn_data_out_rsci_d_207 , chn_data_out_rsci_d_206 , chn_data_out_rsci_d_205_202
      , chn_data_out_rsci_d_201_199 , chn_data_out_rsci_d_198_193 , chn_data_out_rsci_d_192
      , chn_data_out_rsci_d_191 , chn_data_out_rsci_d_190 , chn_data_out_rsci_d_189_186
      , chn_data_out_rsci_d_185_183 , chn_data_out_rsci_d_182_177 , chn_data_out_rsci_d_176
      , chn_data_out_rsci_d_175 , chn_data_out_rsci_d_174 , chn_data_out_rsci_d_173_170
      , chn_data_out_rsci_d_169_167 , chn_data_out_rsci_d_166_161 , chn_data_out_rsci_d_160
      , chn_data_out_rsci_d_159 , chn_data_out_rsci_d_158 , chn_data_out_rsci_d_157_154
      , chn_data_out_rsci_d_153_151 , chn_data_out_rsci_d_150_145 , chn_data_out_rsci_d_144
      , chn_data_out_rsci_d_143 , chn_data_out_rsci_d_142 , chn_data_out_rsci_d_141_138
      , chn_data_out_rsci_d_137_135 , chn_data_out_rsci_d_134_129 , chn_data_out_rsci_d_128
      , chn_data_out_rsci_d_127 , chn_data_out_rsci_d_126 , chn_data_out_rsci_d_125_122
      , chn_data_out_rsci_d_121_119 , chn_data_out_rsci_d_118_113 , chn_data_out_rsci_d_112
      , chn_data_out_rsci_d_111 , chn_data_out_rsci_d_110 , chn_data_out_rsci_d_109_106
      , chn_data_out_rsci_d_105_103 , chn_data_out_rsci_d_102_97 , chn_data_out_rsci_d_96
      , chn_data_out_rsci_d_95 , chn_data_out_rsci_d_94 , chn_data_out_rsci_d_93_90
      , chn_data_out_rsci_d_89_87 , chn_data_out_rsci_d_86_81 , chn_data_out_rsci_d_80
      , chn_data_out_rsci_d_79 , chn_data_out_rsci_d_78 , chn_data_out_rsci_d_77_74
      , chn_data_out_rsci_d_73_71 , chn_data_out_rsci_d_70_65 , chn_data_out_rsci_d_64
      , chn_data_out_rsci_d_63 , chn_data_out_rsci_d_62 , chn_data_out_rsci_d_61_58
      , chn_data_out_rsci_d_57_55 , chn_data_out_rsci_d_54_49 , chn_data_out_rsci_d_48
      , chn_data_out_rsci_d_47 , chn_data_out_rsci_d_46 , chn_data_out_rsci_d_45_42
      , chn_data_out_rsci_d_41_39 , chn_data_out_rsci_d_38_33 , chn_data_out_rsci_d_32
      , chn_data_out_rsci_d_31 , chn_data_out_rsci_d_30 , chn_data_out_rsci_d_29_26
      , chn_data_out_rsci_d_25_23 , chn_data_out_rsci_d_22_17 , chn_data_out_rsci_d_16
      , chn_data_out_rsci_d_15 , chn_data_out_rsci_d_14 , chn_data_out_rsci_d_13_10
      , chn_data_out_rsci_d_9_7 , chn_data_out_rsci_d_6_1 , chn_data_out_rsci_d_0};
  CSC_mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd2)) cfg_truncate_rsci (
      .d(cfg_truncate_rsci_d),
      .z(cfg_truncate_rsc_z)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg
      (
      .a(nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg (
      .a(nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg
      (
      .a(nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg (
      .a(nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg
      (
      .a(nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg (
      .a(nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg (
      .a(nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_a_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg (
      .a(nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_4_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_b_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg
      (
      .a(nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s[4:0]),
      .z(m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg (
      .a(nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_a_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg (
      .a(nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_3_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_b_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg
      (
      .a(nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s[4:0]),
      .z(m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg (
      .a(nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_a_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg (
      .a(nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_2_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_b_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg
      (
      .a(nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s[4:0]),
      .z(m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg (
      .a(nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_a_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg (
      .a(nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row3_1_FpAdd_6U_10U_3_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_3_b_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg (
      .a(nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_a_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg (
      .a(nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_4_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_b_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg (
      .a(nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_a_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg (
      .a(nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_3_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_b_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg (
      .a(nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_a_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg (
      .a(nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_2_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_b_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg (
      .a(nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_a_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg (
      .a(nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row2_1_FpAdd_6U_10U_2_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_2_b_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_a_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_b_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_a_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_b_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_a_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_b_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_a_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row1_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_1_b_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_a_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_b_int_mant_p1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_a_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_b_int_mant_p1_3_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_a_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_b_int_mant_p1_2_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_a_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_m_row0_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_b_int_mant_p1_1_sva_mx0w0)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg
      (
      .a(nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg (
      .a(nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_l #(.width_a(32'sd9),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd10)) m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg
      (
      .a(nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_a[8:0]),
      .s(nl_m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_rg_s[4:0]),
      .z(m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_16_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_16_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_15_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_15_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_14_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_14_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_13_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_13_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_12_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_12_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_11_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_11_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_10_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_10_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_9_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_9_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_8_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_8_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_7_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_7_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_6_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_6_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_5_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_5_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_4_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_4_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_3_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_3_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_2_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_2_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0)
    );
  CSC_mgc_shift_r #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_s(32'sd2),
  .width_z(32'sd21)) data_truncate_1_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg
      (
      .a(nl_data_truncate_1_IntShiftRight_18U_2U_16U_mbits_fixed_rshift_rg_a[20:0]),
      .s(cfg_truncate_rsci_d),
      .z(IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0)
    );
  CSC_leading_sign_10_0  m_row0_1_leading_sign_10_0_rg (
      .mantissa(nl_m_row0_1_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_32)
    );
  CSC_leading_sign_10_0  m_row0_1_leading_sign_10_0_1_rg (
      .mantissa(nl_m_row0_1_leading_sign_10_0_1_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_33)
    );
  CSC_leading_sign_10_0  m_row0_2_leading_sign_10_0_rg (
      .mantissa(nl_m_row0_2_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_34)
    );
  CSC_leading_sign_10_0  m_row0_2_leading_sign_10_0_1_rg (
      .mantissa(nl_m_row0_2_leading_sign_10_0_1_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_35)
    );
  CSC_leading_sign_10_0  m_row0_3_leading_sign_10_0_rg (
      .mantissa(nl_m_row0_3_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_36)
    );
  CSC_leading_sign_10_0  m_row0_3_leading_sign_10_0_1_rg (
      .mantissa(nl_m_row0_3_leading_sign_10_0_1_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_37)
    );
  CSC_leading_sign_10_0  m_row0_4_leading_sign_10_0_rg (
      .mantissa(nl_m_row0_4_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_38)
    );
  CSC_leading_sign_10_0  m_row0_4_leading_sign_10_0_1_rg (
      .mantissa(nl_m_row0_4_leading_sign_10_0_1_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_39)
    );
  CSC_leading_sign_10_0  m_row1_1_leading_sign_10_0_2_rg (
      .mantissa(nl_m_row1_1_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_40)
    );
  CSC_leading_sign_10_0  m_row1_2_leading_sign_10_0_2_rg (
      .mantissa(nl_m_row1_2_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_41)
    );
  CSC_leading_sign_10_0  m_row1_3_leading_sign_10_0_2_rg (
      .mantissa(nl_m_row1_3_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_42)
    );
  CSC_leading_sign_10_0  m_row1_4_leading_sign_10_0_2_rg (
      .mantissa(nl_m_row1_4_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_43)
    );
  CSC_leading_sign_10_0  m_row3_1_leading_sign_10_0_7_rg (
      .mantissa(nl_m_row3_1_leading_sign_10_0_7_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_44)
    );
  CSC_leading_sign_10_0  m_row3_2_leading_sign_10_0_7_rg (
      .mantissa(nl_m_row3_2_leading_sign_10_0_7_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_45)
    );
  CSC_leading_sign_10_0  m_row3_3_leading_sign_10_0_7_rg (
      .mantissa(nl_m_row3_3_leading_sign_10_0_7_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_46)
    );
  CSC_leading_sign_10_0  m_row3_4_leading_sign_10_0_7_rg (
      .mantissa(nl_m_row3_4_leading_sign_10_0_7_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_47)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row0_1_FpNormalize_6U_23U_else_lshift_rg (
      .a(FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_32),
      .z(m_row0_1_FpNormalize_6U_23U_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row0_1_leading_sign_23_0_rg (
      .mantissa(FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_32)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row0_2_FpNormalize_6U_23U_else_lshift_rg (
      .a(FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_33),
      .z(m_row0_2_FpNormalize_6U_23U_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row0_2_leading_sign_23_0_rg (
      .mantissa(FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_33)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row0_3_FpNormalize_6U_23U_else_lshift_rg (
      .a(FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_34),
      .z(m_row0_3_FpNormalize_6U_23U_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row0_3_leading_sign_23_0_rg (
      .mantissa(FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_34)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row0_4_FpNormalize_6U_23U_else_lshift_rg (
      .a(FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_35),
      .z(m_row0_4_FpNormalize_6U_23U_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row0_4_leading_sign_23_0_rg (
      .mantissa(FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_35)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row1_1_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_36),
      .z(m_row1_1_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row1_1_leading_sign_23_0_1_rg (
      .mantissa(FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_36)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row1_2_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_37),
      .z(m_row1_2_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row1_2_leading_sign_23_0_1_rg (
      .mantissa(FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_37)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row1_3_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_38),
      .z(m_row1_3_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row1_3_leading_sign_23_0_1_rg (
      .mantissa(FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_38)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row1_4_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_39),
      .z(m_row1_4_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row1_4_leading_sign_23_0_1_rg (
      .mantissa(FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_39)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row2_1_FpNormalize_6U_23U_2_else_lshift_rg (
      .a(FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_40),
      .z(m_row2_1_FpNormalize_6U_23U_2_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row2_1_leading_sign_23_0_2_rg (
      .mantissa(FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_40)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row2_2_FpNormalize_6U_23U_2_else_lshift_rg (
      .a(FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_41),
      .z(m_row2_2_FpNormalize_6U_23U_2_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row2_2_leading_sign_23_0_2_rg (
      .mantissa(FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_41)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row2_3_FpNormalize_6U_23U_2_else_lshift_rg (
      .a(FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_42),
      .z(m_row2_3_FpNormalize_6U_23U_2_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row2_3_leading_sign_23_0_2_rg (
      .mantissa(FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_42)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row2_4_FpNormalize_6U_23U_2_else_lshift_rg (
      .a(FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_43),
      .z(m_row2_4_FpNormalize_6U_23U_2_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row2_4_leading_sign_23_0_2_rg (
      .mantissa(FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_43)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row3_1_FpNormalize_6U_23U_3_else_lshift_rg (
      .a(FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_44),
      .z(m_row3_1_FpNormalize_6U_23U_3_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row3_1_leading_sign_23_0_3_rg (
      .mantissa(FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_44)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row3_2_FpNormalize_6U_23U_3_else_lshift_rg (
      .a(FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_45),
      .z(m_row3_2_FpNormalize_6U_23U_3_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row3_2_leading_sign_23_0_3_rg (
      .mantissa(FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_45)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row3_3_FpNormalize_6U_23U_3_else_lshift_rg (
      .a(FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_46),
      .z(m_row3_3_FpNormalize_6U_23U_3_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row3_3_leading_sign_23_0_3_rg (
      .mantissa(FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_46)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) m_row3_4_FpNormalize_6U_23U_3_else_lshift_rg (
      .a(FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_47),
      .z(m_row3_4_FpNormalize_6U_23U_3_else_lshift_itm)
    );
  CSC_leading_sign_23_0  m_row3_4_leading_sign_23_0_3_rg (
      .mantissa(FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_47)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col0_1_FpNormalize_6U_23U_4_else_lshift_rg (
      .a(nl_o_col0_1_FpNormalize_6U_23U_4_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_48),
      .z(o_col0_1_FpNormalize_6U_23U_4_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col0_1_leading_sign_23_0_4_rg (
      .mantissa(nl_o_col0_1_leading_sign_23_0_4_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_48)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col0_2_FpNormalize_6U_23U_4_else_lshift_rg (
      .a(nl_o_col0_2_FpNormalize_6U_23U_4_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_49),
      .z(o_col0_2_FpNormalize_6U_23U_4_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col0_2_leading_sign_23_0_4_rg (
      .mantissa(nl_o_col0_2_leading_sign_23_0_4_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_49)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col0_3_FpNormalize_6U_23U_4_else_lshift_rg (
      .a(nl_o_col0_3_FpNormalize_6U_23U_4_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_50),
      .z(o_col0_3_FpNormalize_6U_23U_4_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col0_3_leading_sign_23_0_4_rg (
      .mantissa(nl_o_col0_3_leading_sign_23_0_4_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_50)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col0_4_FpNormalize_6U_23U_4_else_lshift_rg (
      .a(nl_o_col0_4_FpNormalize_6U_23U_4_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_51),
      .z(o_col0_4_FpNormalize_6U_23U_4_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col0_4_leading_sign_23_0_4_rg (
      .mantissa(nl_o_col0_4_leading_sign_23_0_4_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_51)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col1_1_FpNormalize_6U_23U_5_else_lshift_rg (
      .a(nl_o_col1_1_FpNormalize_6U_23U_5_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_52),
      .z(o_col1_1_FpNormalize_6U_23U_5_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col1_1_leading_sign_23_0_5_rg (
      .mantissa(nl_o_col1_1_leading_sign_23_0_5_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_52)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col1_2_FpNormalize_6U_23U_5_else_lshift_rg (
      .a(nl_o_col1_2_FpNormalize_6U_23U_5_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_53),
      .z(o_col1_2_FpNormalize_6U_23U_5_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col1_2_leading_sign_23_0_5_rg (
      .mantissa(nl_o_col1_2_leading_sign_23_0_5_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_53)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col1_3_FpNormalize_6U_23U_5_else_lshift_rg (
      .a(nl_o_col1_3_FpNormalize_6U_23U_5_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_54),
      .z(o_col1_3_FpNormalize_6U_23U_5_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col1_3_leading_sign_23_0_5_rg (
      .mantissa(nl_o_col1_3_leading_sign_23_0_5_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_54)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col1_4_FpNormalize_6U_23U_5_else_lshift_rg (
      .a(nl_o_col1_4_FpNormalize_6U_23U_5_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_55),
      .z(o_col1_4_FpNormalize_6U_23U_5_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col1_4_leading_sign_23_0_5_rg (
      .mantissa(nl_o_col1_4_leading_sign_23_0_5_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_55)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col2_1_FpNormalize_6U_23U_6_else_lshift_rg (
      .a(nl_o_col2_1_FpNormalize_6U_23U_6_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_56),
      .z(o_col2_1_FpNormalize_6U_23U_6_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col2_1_leading_sign_23_0_6_rg (
      .mantissa(nl_o_col2_1_leading_sign_23_0_6_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_56)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col2_2_FpNormalize_6U_23U_6_else_lshift_rg (
      .a(nl_o_col2_2_FpNormalize_6U_23U_6_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_57),
      .z(o_col2_2_FpNormalize_6U_23U_6_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col2_2_leading_sign_23_0_6_rg (
      .mantissa(nl_o_col2_2_leading_sign_23_0_6_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_57)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col2_3_FpNormalize_6U_23U_6_else_lshift_rg (
      .a(nl_o_col2_3_FpNormalize_6U_23U_6_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_58),
      .z(o_col2_3_FpNormalize_6U_23U_6_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col2_3_leading_sign_23_0_6_rg (
      .mantissa(nl_o_col2_3_leading_sign_23_0_6_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_58)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col2_4_FpNormalize_6U_23U_6_else_lshift_rg (
      .a(nl_o_col2_4_FpNormalize_6U_23U_6_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_59),
      .z(o_col2_4_FpNormalize_6U_23U_6_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col2_4_leading_sign_23_0_6_rg (
      .mantissa(nl_o_col2_4_leading_sign_23_0_6_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_59)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col3_1_FpNormalize_6U_23U_7_else_lshift_rg (
      .a(nl_o_col3_1_FpNormalize_6U_23U_7_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_60),
      .z(o_col3_1_FpNormalize_6U_23U_7_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col3_1_leading_sign_23_0_7_rg (
      .mantissa(nl_o_col3_1_leading_sign_23_0_7_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_60)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col3_2_FpNormalize_6U_23U_7_else_lshift_rg (
      .a(nl_o_col3_2_FpNormalize_6U_23U_7_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_61),
      .z(o_col3_2_FpNormalize_6U_23U_7_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col3_2_leading_sign_23_0_7_rg (
      .mantissa(nl_o_col3_2_leading_sign_23_0_7_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_61)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col3_3_FpNormalize_6U_23U_7_else_lshift_rg (
      .a(nl_o_col3_3_FpNormalize_6U_23U_7_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_62),
      .z(o_col3_3_FpNormalize_6U_23U_7_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col3_3_leading_sign_23_0_7_rg (
      .mantissa(nl_o_col3_3_leading_sign_23_0_7_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_62)
    );
  CSC_mgc_shift_l #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) o_col3_4_FpNormalize_6U_23U_7_else_lshift_rg (
      .a(nl_o_col3_4_FpNormalize_6U_23U_7_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_63),
      .z(o_col3_4_FpNormalize_6U_23U_7_else_lshift_itm)
    );
  CSC_leading_sign_23_0  o_col3_4_leading_sign_23_0_7_rg (
      .mantissa(nl_o_col3_4_leading_sign_23_0_7_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_63)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_1_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_1_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_1_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_1_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_1_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_2_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_2_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_2_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_2_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_2_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_3_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_3_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_3_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_3_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_3_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_4_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_4_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_4_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_4_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_4_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_5_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_5_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_5_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_5_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_5_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_6_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_6_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_6_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_6_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_6_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_7_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_7_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_7_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_7_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_7_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_8_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_8_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_8_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_8_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_8_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_9_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_9_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_9_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_9_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_9_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_10_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_10_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_10_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_10_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_10_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_11_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_11_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_11_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_11_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_11_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_12_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_12_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_12_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_12_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_12_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_13_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_13_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_13_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_13_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_13_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_14_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_14_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_14_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_14_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_14_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_15_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_15_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_15_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_15_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_15_sva)
    );
  CSC_mgc_shift_r #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg
      (
      .a(nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_a[10:0]),
      .s(nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd11)) data_truncate_16_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_guard_mask_sva)
    );
  CSC_mgc_shift_l #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) data_truncate_16_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_data_truncate_16_FpMantDecShiftRight_10U_6U_10U_least_mask_lshift_rg_s[3:0]),
      .z(FpMantDecShiftRight_10U_6U_10U_least_mask_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg (
      .a(nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_1_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_addend_larger_asn_19_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg (
      .a(nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_1_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_a_int_mant_p1_1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg (
      .a(nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_2_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_addend_larger_asn_13_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg (
      .a(nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_2_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_a_int_mant_p1_2_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg (
      .a(nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_3_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_addend_larger_asn_7_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg (
      .a(nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_3_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_a_int_mant_p1_3_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg (
      .a(nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_4_FpAdd_6U_10U_4_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_addend_larger_asn_1_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg (
      .a(nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col0_4_FpAdd_6U_10U_4_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_4_a_int_mant_p1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg (
      .a(nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_1_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_addend_larger_asn_19_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg (
      .a(nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_1_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_a_int_mant_p1_1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg (
      .a(nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_2_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_addend_larger_asn_13_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg (
      .a(nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_2_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_a_int_mant_p1_2_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg (
      .a(nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_3_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_addend_larger_asn_7_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg (
      .a(nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_3_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_a_int_mant_p1_3_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg (
      .a(nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_4_FpAdd_6U_10U_5_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_addend_larger_asn_1_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg (
      .a(nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col1_4_FpAdd_6U_10U_5_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_5_a_int_mant_p1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg (
      .a(nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_1_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_addend_larger_asn_19_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg (
      .a(nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_1_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_a_int_mant_p1_1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg (
      .a(nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_2_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_addend_larger_asn_13_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg (
      .a(nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_2_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_a_int_mant_p1_2_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg (
      .a(nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_3_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_addend_larger_asn_7_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg (
      .a(nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_3_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_a_int_mant_p1_3_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg (
      .a(nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_4_FpAdd_6U_10U_6_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_addend_larger_asn_1_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg (
      .a(nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col2_4_FpAdd_6U_10U_6_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_6_a_int_mant_p1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg (
      .a(nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_1_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_addend_larger_asn_19_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg (
      .a(nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_1_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_a_int_mant_p1_1_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg (
      .a(nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_2_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_addend_larger_asn_13_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg (
      .a(nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_2_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_a_int_mant_p1_2_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg (
      .a(nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_3_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_addend_larger_asn_7_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg (
      .a(nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_3_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_a_int_mant_p1_3_sva)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg (
      .a(nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_4_FpAdd_6U_10U_7_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_addend_larger_asn_1_mx0w1)
    );
  CSC_mgc_shift_bl #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg (
      .a(nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_o_col3_4_FpAdd_6U_10U_7_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(FpAdd_6U_10U_7_a_int_mant_p1_sva)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci NV_NVDLA_CSC_pra_cell_core_chn_data_in_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_in_rsc_z(chn_data_in_rsc_z),
      .chn_data_in_rsc_vz(chn_data_in_rsc_vz),
      .chn_data_in_rsc_lz(chn_data_in_rsc_lz),
      .chn_data_in_rsci_oswt(chn_data_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_data_in_rsci_iswt0(chn_data_in_rsci_iswt0),
      .chn_data_in_rsci_bawt(chn_data_in_rsci_bawt),
      .chn_data_in_rsci_wen_comp(chn_data_in_rsci_wen_comp),
      .chn_data_in_rsci_ld_core_psct(chn_data_in_rsci_ld_core_psct),
      .chn_data_in_rsci_d_mxwt(chn_data_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_out_rsc_z(chn_data_out_rsc_z),
      .chn_data_out_rsc_vz(chn_data_out_rsc_vz),
      .chn_data_out_rsc_lz(chn_data_out_rsc_lz),
      .chn_data_out_rsci_oswt(chn_data_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_data_out_rsci_iswt0(chn_data_out_rsci_iswt0),
      .chn_data_out_rsci_bawt(chn_data_out_rsci_bawt),
      .chn_data_out_rsci_wen_comp(chn_data_out_rsci_wen_comp),
      .chn_data_out_rsci_ld_core_psct(reg_chn_data_out_rsci_ld_core_psct_cse),
      .chn_data_out_rsci_d(nl_NV_NVDLA_CSC_pra_cell_core_chn_data_out_rsci_inst_chn_data_out_rsci_d[255:0])
    );
  NV_NVDLA_CSC_pra_cell_core_staller NV_NVDLA_CSC_pra_cell_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_data_in_rsci_wen_comp(chn_data_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_data_out_rsci_wen_comp(chn_data_out_rsci_wen_comp)
    );
  NV_NVDLA_CSC_pra_cell_core_core_fsm NV_NVDLA_CSC_pra_cell_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_16 = and_dcpl_3 & (~ data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1)
      & data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva)
      , (FpAdd_6U_10U_4_o_expo_1_lpi_2[0])}) + 5'b1)), and_16);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb } @rose(nvdla_core_clk);
  assign and_19 = and_dcpl_3 & data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_1 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva)
      , (FpAdd_6U_10U_5_o_expo_1_lpi_2[0])}) + 5'b1)), and_19);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_1 } @rose(nvdla_core_clk);
  assign and_22 = and_dcpl_3 & data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_2 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva)
      , (FpAdd_6U_10U_6_o_expo_1_lpi_2[0])}) + 5'b1)), and_22);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_2 } @rose(nvdla_core_clk);
  assign and_25 = and_dcpl_3 & data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_3 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva)
      , (FpAdd_6U_10U_7_o_expo_1_lpi_2[0])}) + 5'b1)), and_25);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_3 } @rose(nvdla_core_clk);
  assign and_28 = and_dcpl_3 & data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_4 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva)
      , (FpAdd_6U_10U_4_o_expo_2_lpi_2[0])}) + 5'b1)), and_28);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_5_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_4 } @rose(nvdla_core_clk);
  assign and_31 = and_dcpl_3 & data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_5 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva)
      , (FpAdd_6U_10U_5_o_expo_2_lpi_2[0])}) + 5'b1)), and_31);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_6_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_5 } @rose(nvdla_core_clk);
  assign and_34 = and_dcpl_3 & data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_6 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva)
      , (FpAdd_6U_10U_6_o_expo_2_lpi_2[0])}) + 5'b1)), and_34);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_7_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_6 } @rose(nvdla_core_clk);
  assign and_37 = and_dcpl_3 & data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_7 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva)
      , (FpAdd_6U_10U_7_o_expo_2_lpi_2[0])}) + 5'b1)), and_37);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_8_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_7 } @rose(nvdla_core_clk);
  assign and_40 = and_dcpl_3 & data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_8 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva)
      , (FpAdd_6U_10U_4_o_expo_3_lpi_2[0])}) + 5'b1)), and_40);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_9_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_8 } @rose(nvdla_core_clk);
  assign and_43 = and_dcpl_3 & (~ data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_9 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva)
      , (FpAdd_6U_10U_5_o_expo_3_lpi_2[0])}) + 5'b1)), and_43);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_10_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_9 } @rose(nvdla_core_clk);
  assign and_46 = and_dcpl_3 & data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1)
      & (~ data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1);
  assign shift_0_prb_10 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva)
      , (FpAdd_6U_10U_6_o_expo_3_lpi_2[0])}) + 5'b1)), and_46);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_11_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_10 } @rose(nvdla_core_clk);
  assign and_49 = and_dcpl_3 & (~(data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1
      | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1)) & data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign shift_0_prb_11 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva)
      , (FpAdd_6U_10U_7_o_expo_3_lpi_2[0])}) + 5'b1)), and_49);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_12_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_11 } @rose(nvdla_core_clk);
  assign and_52 = and_dcpl_3 & data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_12 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva)
      , (FpAdd_6U_10U_4_o_expo_lpi_2[0])}) + 5'b1)), and_52);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_13_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_12 } @rose(nvdla_core_clk);
  assign and_55 = and_dcpl_3 & data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_13 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva)
      , (FpAdd_6U_10U_5_o_expo_lpi_2[0])}) + 5'b1)), and_55);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_14_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_13 } @rose(nvdla_core_clk);
  assign and_58 = and_dcpl_3 & data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_14 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva)
      , (FpAdd_6U_10U_6_o_expo_lpi_2[0])}) + 5'b1)), and_58);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_15_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_14 } @rose(nvdla_core_clk);
  assign and_61 = and_dcpl_3 & data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & (~ data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1) &
      (~ data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign shift_0_prb_15 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva)
      , (FpAdd_6U_10U_7_o_expo_lpi_2[0])}) + 5'b1)), and_61);
  // assert(shift > 0) - ../include/nvdla_float.h: line 340
  // PSL data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln340_assert_shift_gt_0 : assert { shift_0_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_2 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_2 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_3 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_4 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_4 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_5 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_6 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_6 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_7 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row0_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_8 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_8 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_9 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_10 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_10 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_11 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_12 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_12 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_13 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_14 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_14 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_15 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row1_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_16 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_16 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_17 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_17 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_18 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_18 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_19 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_19 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_20 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_20 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_21 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_21 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_22 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_22 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_23 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row2_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_24 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_6 : assert { iExpoWidth_oExpoWidth_prb_24 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_25 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7 : assert { iExpoWidth_oExpoWidth_prb_25 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_26 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_6 : assert { iExpoWidth_oExpoWidth_prb_26 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_27 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7 : assert { iExpoWidth_oExpoWidth_prb_27 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_28 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_6 : assert { iExpoWidth_oExpoWidth_prb_28 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_29 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7 : assert { iExpoWidth_oExpoWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_30 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_6 : assert { iExpoWidth_oExpoWidth_prb_30 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_31 = m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1;
  // assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 477
  // PSL m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7 : assert { iExpoWidth_oExpoWidth_prb_31 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row0_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_1 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row0_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_1 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_2 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row0_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_2 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_3 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row0_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_3 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_4 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL m_row1_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_4 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_5 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL m_row1_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_5 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_6 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL m_row1_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_6 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_7 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL m_row1_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb_7 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_8 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row2_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_8 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_9 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row2_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_9 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_10 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row2_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_10 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_11 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row2_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_11 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_12 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row3_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_12 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_13 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row3_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_13 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_14 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row3_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_14 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_15 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_15 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_16 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col0_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_16 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_17 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col0_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_17 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_18 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col0_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_18 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_19 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col0_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_19 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_20 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL o_col1_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_20 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_21 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL o_col1_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_21 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_22 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL o_col1_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_22 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_23 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 257
  // PSL o_col1_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln257_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_23 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_24 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col2_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_4 : assert { oWidth_mWidth_prb_24 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_25 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col2_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_4 : assert { oWidth_mWidth_prb_25 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_26 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col2_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_4 : assert { oWidth_mWidth_prb_26 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_27 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col2_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_4 : assert { oWidth_mWidth_prb_27 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_28 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col3_1_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5 : assert { oWidth_mWidth_prb_28 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_29 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col3_2_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5 : assert { oWidth_mWidth_prb_29 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_30 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col3_3_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5 : assert { oWidth_mWidth_prb_30 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_31 = o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1;
  // assert(oWidth > mWidth) - ../include/nvdla_int.h: line 274
  // PSL o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5 : assert { oWidth_mWidth_prb_31 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_32 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_1_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_32 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_33 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_2_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_33 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_34 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_3_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_34 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_35 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_35 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_36 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_5_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_36 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_37 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_6_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_37 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_38 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_7_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_38 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_39 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_8_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_39 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_40 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_9_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_40 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_41 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_10_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_41 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_42 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_11_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_42 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_43 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_12_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_43 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_44 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_13_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_44 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_45 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_14_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_45 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_46 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_15_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_46 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_47 = data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1;
  // assert(iExpoWidth > oExpoWidth) - ../include/nvdla_float.h: line 630
  // PSL data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_47 } @rose(nvdla_core_clk);
  assign chn_data_out_and_cse = core_wen & (~(and_dcpl_64 | (~ main_stage_v_4)));
  assign FpAdd_6U_10U_and_cse = core_wen & (~ and_dcpl_64) & mux_tmp_49;
  assign and_358_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp;
  assign and_360_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp);
  assign nor_57_cse = ~((cfg_precision!=2'b10));
  assign or_99_cse = IsNaN_6U_10U_1_land_1_lpi_1_dfm | IsNaN_6U_10U_land_1_lpi_1_dfm;
  assign and_370_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_79;
  assign and_374_rgt = and_dcpl_90 & and_dcpl_88 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_tmp);
  assign and_383_rgt = and_dcpl_99 & and_dcpl_94 & and_dcpl_92;
  assign and_386_rgt = and_dcpl_102 & and_dcpl_101;
  assign and_388_rgt = or_dcpl_70 & or_181_cse;
  assign and_390_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp;
  assign and_392_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp);
  assign or_109_cse = IsNaN_6U_10U_1_land_2_lpi_1_dfm | IsNaN_6U_10U_land_2_lpi_1_dfm;
  assign and_401_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_110;
  assign and_404_rgt = and_dcpl_120 & and_dcpl_88 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp);
  assign and_413_rgt = and_dcpl_129 & and_dcpl_124 & and_dcpl_122;
  assign and_416_rgt = and_dcpl_132 & and_dcpl_88 & IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
  assign and_418_rgt = (or_dcpl_1 | IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp) & or_181_cse;
  assign and_420_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp;
  assign and_422_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp);
  assign or_119_cse = IsNaN_6U_10U_1_land_3_lpi_1_dfm | IsNaN_6U_10U_land_3_lpi_1_dfm;
  assign and_431_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_140;
  assign and_434_rgt = and_dcpl_150 & and_dcpl_88 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp);
  assign and_443_rgt = and_dcpl_159 & and_dcpl_154 & and_dcpl_152;
  assign and_446_rgt = and_dcpl_162 & and_dcpl_161;
  assign and_448_rgt = or_dcpl_92 & or_181_cse;
  assign and_450_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp;
  assign and_452_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp);
  assign and_454_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp;
  assign and_456_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp);
  assign and_459_rgt = or_dcpl_93 & or_181_cse;
  assign and_461_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp;
  assign and_463_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp);
  assign and_466_rgt = or_dcpl_94 & or_181_cse;
  assign and_468_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp;
  assign and_470_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp);
  assign and_473_rgt = or_dcpl_95 & or_181_cse;
  assign and_475_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp;
  assign and_477_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp);
  assign and_479_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp;
  assign and_481_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp);
  assign and_484_rgt = (or_dcpl_1 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp) & or_181_cse;
  assign and_486_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp;
  assign and_488_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp);
  assign and_491_rgt = (or_dcpl_1 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp) & or_181_cse;
  assign and_493_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp;
  assign and_495_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp);
  assign and_498_rgt = (or_dcpl_1 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp) & or_181_cse;
  assign and_500_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp;
  assign and_502_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp);
  assign and_504_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp;
  assign and_506_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp);
  assign and_509_rgt = or_dcpl_99 & or_181_cse;
  assign and_511_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp;
  assign and_513_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp);
  assign and_516_rgt = or_dcpl_100 & or_181_cse;
  assign and_518_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp;
  assign and_520_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp);
  assign and_523_rgt = (or_dcpl_1 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp) & or_181_cse;
  assign and_525_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp;
  assign and_527_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp);
  assign IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse = and_dcpl_245 | and_dcpl_78;
  assign IsNaN_6U_10U_6_aelse_and_8_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & mux_tmp_49;
  assign nor_546_cse = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ main_stage_v_1));
  assign or_nl = main_stage_v_1 | or_181_cse;
  assign mux_67_cse = MUX_s_1_2_2(nor_546_cse, (or_nl), chn_data_in_rsci_bawt);
  assign FpAdd_6U_10U_3_a_int_mant_p1_and_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & mux_67_cse;
  assign nor_70_cse = ~(IsNaN_6U_10U_6_land_3_lpi_1_dfm | (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm));
  assign or_134_cse = nor_70_cse | IsNaN_6U_10U_6_land_3_lpi_1_dfm;
  assign and_537_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_246;
  assign and_540_rgt = and_dcpl_256 & and_dcpl_88 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign and_548_rgt = and_dcpl_264 & and_dcpl_259 & and_dcpl_238;
  assign and_551_rgt = and_dcpl_267 & and_dcpl_88 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_cse = core_wen & (and_dcpl_269
      | and_dcpl_270 | and_dcpl_271) & mux_tmp_76;
  assign mux_79_cse = MUX_s_1_2_2(main_stage_v_1, chn_data_in_rsci_bawt, or_181_cse);
  assign FpAdd_6U_10U_3_a_int_mant_p1_and_7_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & mux_79_cse;
  assign or_152_cse = IsNaN_6U_10U_7_land_2_lpi_1_dfm | IsNaN_6U_10U_6_land_2_lpi_1_dfm;
  assign and_564_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_272;
  assign and_567_rgt = and_dcpl_282 & and_dcpl_281;
  assign and_575_rgt = and_dcpl_290 & and_dcpl_285 & and_dcpl_231;
  assign and_578_rgt = and_dcpl_293 & and_dcpl_88 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_3_cse = core_wen & (and_dcpl_295
      | and_dcpl_296 | and_dcpl_297) & mux_tmp_88;
  assign nor_82_cse = ~(IsNaN_6U_10U_6_land_1_lpi_1_dfm | (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm));
  assign and_590_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_298;
  assign and_593_rgt = and_dcpl_308 & and_dcpl_307;
  assign and_601_rgt = and_dcpl_316 & and_dcpl_311 & and_dcpl_224;
  assign and_604_rgt = and_dcpl_319 & and_dcpl_88 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_6_cse = core_wen & (and_dcpl_321
      | and_dcpl_322 | and_dcpl_323) & mux_tmp_100;
  assign or_181_cse = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt;
  assign or_183_cse = IsNaN_6U_10U_5_land_3_lpi_1_dfm | IsNaN_6U_10U_4_land_3_lpi_1_dfm;
  assign and_610_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_324;
  assign and_612_rgt = and_dcpl_150 & and_dcpl_88 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign and_614_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_213;
  assign and_616_rgt = and_dcpl_256 & and_dcpl_88 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp);
  assign or_1963_cse = IsNaN_6U_10U_5_land_3_lpi_1_dfm_3 | IsNaN_6U_10U_4_land_3_lpi_1_dfm_3;
  assign and_2591_cse = or_1963_cse & main_stage_v_1;
  assign mux_109_nl = MUX_s_1_2_2(not_tmp_109, or_tmp_170, or_tmp_39);
  assign mux_110_nl = MUX_s_1_2_2(not_tmp_109, or_tmp_170, or_183_cse);
  assign mux_111_nl = MUX_s_1_2_2((mux_110_nl), (mux_109_nl), nor_57_cse);
  assign mux_112_nl = MUX_s_1_2_2(not_tmp_109, (mux_111_nl), chn_data_in_rsci_bawt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_cse = core_wen & (and_dcpl_333
      | and_dcpl_78 | and_dcpl_214) & (mux_112_nl);
  assign or_196_cse = IsNaN_6U_10U_5_land_2_lpi_1_dfm | IsNaN_6U_10U_4_land_2_lpi_1_dfm;
  assign and_620_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_334;
  assign and_622_rgt = and_dcpl_120 & and_dcpl_88 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
  assign and_624_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_206;
  assign and_626_rgt = and_dcpl_282 & and_dcpl_88 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign or_1962_cse = IsNaN_6U_10U_5_land_2_lpi_1_dfm_3 | IsNaN_6U_10U_4_land_2_lpi_1_dfm_3;
  assign and_2588_cse = or_1962_cse & main_stage_v_1;
  assign mux_118_nl = MUX_s_1_2_2(not_tmp_112, or_tmp_183, or_tmp_36);
  assign mux_119_nl = MUX_s_1_2_2(not_tmp_112, or_tmp_183, or_196_cse);
  assign mux_120_nl = MUX_s_1_2_2((mux_119_nl), (mux_118_nl), nor_57_cse);
  assign mux_121_nl = MUX_s_1_2_2(not_tmp_112, (mux_120_nl), chn_data_in_rsci_bawt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_3_cse = core_wen & (and_dcpl_343
      | and_dcpl_78 | and_dcpl_207) & (mux_121_nl);
  assign or_209_cse = IsNaN_6U_10U_5_land_1_lpi_1_dfm | IsNaN_6U_10U_4_land_1_lpi_1_dfm;
  assign and_630_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_344;
  assign and_632_rgt = and_dcpl_90 & and_dcpl_88 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
  assign and_634_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_199;
  assign and_636_rgt = and_dcpl_308 & and_dcpl_88 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp);
  assign or_1961_cse = IsNaN_6U_10U_5_land_1_lpi_1_dfm_3 | IsNaN_6U_10U_4_land_1_lpi_1_dfm_3;
  assign and_2585_cse = or_1961_cse & main_stage_v_1;
  assign mux_127_nl = MUX_s_1_2_2(not_tmp_115, or_tmp_196, or_tmp_33);
  assign mux_128_nl = MUX_s_1_2_2(not_tmp_115, or_tmp_196, or_209_cse);
  assign mux_129_nl = MUX_s_1_2_2((mux_128_nl), (mux_127_nl), nor_57_cse);
  assign mux_130_nl = MUX_s_1_2_2(not_tmp_115, (mux_129_nl), chn_data_in_rsci_bawt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_6_cse = core_wen & (and_dcpl_353
      | and_dcpl_78 | and_dcpl_200) & (mux_130_nl);
  assign or_224_cse = IsNaN_6U_10U_3_land_3_lpi_1_dfm | IsNaN_6U_10U_2_land_3_lpi_1_dfm;
  assign and_640_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_354;
  assign and_642_rgt = and_dcpl_256 & and_dcpl_357;
  assign and_644_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_188;
  assign and_646_rgt = and_dcpl_150 & and_dcpl_88 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign or_1960_cse = IsNaN_6U_10U_3_land_3_lpi_1_dfm_3 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_3;
  assign and_2582_cse = or_1960_cse & main_stage_v_1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse = core_wen & (and_dcpl_363
      | and_dcpl_189 | and_dcpl_364) & mux_tmp_142;
  assign and_649_rgt = and_dcpl_74 & and_dcpl_354;
  assign or_237_cse = IsNaN_6U_10U_3_land_2_lpi_1_dfm | IsNaN_6U_10U_2_land_2_lpi_1_dfm;
  assign and_652_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_366;
  assign and_654_rgt = and_dcpl_282 & and_dcpl_369;
  assign and_656_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_181;
  assign and_658_rgt = and_dcpl_120 & and_dcpl_88 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign or_1959_cse = IsNaN_6U_10U_3_land_2_lpi_1_dfm_3 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_3;
  assign and_2579_cse = or_1959_cse & main_stage_v_1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_3_cse = core_wen & (and_dcpl_375
      | and_dcpl_182 | and_dcpl_376) & mux_tmp_151;
  assign and_661_rgt = and_dcpl_74 & and_dcpl_366;
  assign or_1980_nl = nor_tmp_118 | or_181_cse;
  assign nor_523_nl = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_118));
  assign mux_153_nl = MUX_s_1_2_2((nor_523_nl), (or_1980_nl), chn_data_in_rsci_bawt);
  assign mux_156_nl = MUX_s_1_2_2(mux_67_cse, (mux_153_nl), reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_a_int_mant_p1_and_8_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & (mux_156_nl);
  assign or_256_cse = IsNaN_6U_10U_3_land_1_lpi_1_dfm | IsNaN_6U_10U_2_land_1_lpi_1_dfm;
  assign and_664_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_378;
  assign and_666_rgt = and_dcpl_308 & and_dcpl_381;
  assign and_668_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_174;
  assign and_670_rgt = and_dcpl_90 & and_dcpl_88 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign or_1958_cse = IsNaN_6U_10U_3_land_1_lpi_1_dfm_3 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_3;
  assign and_2576_cse = or_1958_cse & main_stage_v_1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_6_cse = core_wen & (and_dcpl_387
      | and_dcpl_175 | and_dcpl_388) & mux_tmp_162;
  assign and_673_rgt = and_dcpl_74 & and_dcpl_378;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse = core_wen & (((~ mux_tmp_656)
      & or_181_cse) | and_dcpl_391) & mux_tmp_172;
  assign and_676_rgt = and_dcpl_74 & and_dcpl_152;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_3_cse = core_wen & (((~ mux_tmp_657)
      & or_181_cse) | and_dcpl_394) & mux_tmp_179;
  assign and_680_rgt = and_dcpl_74 & and_dcpl_122;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_6_cse = core_wen & (((~ mux_tmp_658)
      & or_181_cse) | and_dcpl_397) & mux_tmp_186;
  assign and_683_rgt = and_dcpl_74 & and_dcpl_92;
  assign and_689_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse);
  assign and_691_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_o_expo_and_cse = core_wen & (~ and_dcpl_64) & mux_468_cse;
  assign and_693_rgt = or_181_cse & (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_3);
  assign and_695_rgt = or_181_cse & (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_3);
  assign and_697_rgt = or_181_cse & (~ IsNaN_6U_10U_4_land_1_lpi_1_dfm_3);
  assign and_699_rgt = or_181_cse & (~ IsNaN_6U_10U_4_land_3_lpi_1_dfm_3);
  assign and_701_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse);
  assign and_703_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse);
  assign and_705_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse);
  assign and_707_rgt = or_181_cse & (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_3);
  assign and_709_rgt = or_181_cse & (~ IsNaN_6U_10U_4_land_2_lpi_1_dfm_3);
  assign and_711_rgt = or_181_cse & (~ reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse);
  assign and_713_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse;
  assign and_715_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse);
  assign and_717_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & IsNaN_6U_10U_2_land_lpi_1_dfm_st_2;
  assign and_719_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_2);
  assign and_721_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & IsNaN_6U_10U_4_land_lpi_1_dfm_st_2;
  assign and_723_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ IsNaN_6U_10U_4_land_lpi_1_dfm_st_2);
  assign and_725_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse;
  assign and_727_rgt = and_dcpl_74 & (~ (cfg_precision[0])) & (~ reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse);
  assign IsNaN_6U_10U_12_aelse_and_4_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & mux_468_cse;
  assign and_733_rgt = and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1;
  assign and_735_rgt = and_dcpl_245 & and_dcpl_449;
  assign FpAdd_6U_10U_4_and_39_ssc = core_wen & (and_733_rgt | and_735_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_737_rgt = and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1;
  assign and_739_rgt = and_dcpl_245 & and_dcpl_453;
  assign FpAdd_6U_10U_4_and_40_ssc = core_wen & (and_737_rgt | and_739_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_741_rgt = and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1;
  assign and_743_rgt = and_dcpl_245 & and_dcpl_457;
  assign FpAdd_6U_10U_4_and_41_ssc = core_wen & (and_741_rgt | and_743_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_745_rgt = and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1;
  assign and_747_rgt = and_dcpl_245 & and_dcpl_461;
  assign FpAdd_6U_10U_4_and_42_ssc = core_wen & (and_745_rgt | and_747_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_749_rgt = and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1;
  assign and_751_rgt = and_dcpl_245 & and_dcpl_465;
  assign FpAdd_6U_10U_5_and_39_ssc = core_wen & (and_749_rgt | and_751_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_753_rgt = and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1;
  assign and_755_rgt = and_dcpl_245 & and_dcpl_469;
  assign FpAdd_6U_10U_5_and_40_ssc = core_wen & (and_753_rgt | and_755_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_757_rgt = and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1;
  assign and_759_rgt = and_dcpl_245 & and_dcpl_473;
  assign FpAdd_6U_10U_5_and_41_ssc = core_wen & (and_757_rgt | and_759_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_761_rgt = and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1;
  assign and_763_rgt = and_dcpl_245 & and_dcpl_477;
  assign FpAdd_6U_10U_5_and_42_ssc = core_wen & (and_761_rgt | and_763_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_765_rgt = and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1;
  assign and_767_rgt = and_dcpl_245 & and_dcpl_481;
  assign FpAdd_6U_10U_6_and_39_ssc = core_wen & (and_765_rgt | and_767_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_769_rgt = and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1;
  assign and_771_rgt = and_dcpl_245 & and_dcpl_485;
  assign FpAdd_6U_10U_6_and_40_ssc = core_wen & (and_769_rgt | and_771_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_773_rgt = and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1;
  assign and_775_rgt = and_dcpl_245 & and_dcpl_489;
  assign FpAdd_6U_10U_6_and_41_ssc = core_wen & (and_773_rgt | and_775_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_777_rgt = and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1;
  assign and_779_rgt = and_dcpl_245 & and_dcpl_493;
  assign FpAdd_6U_10U_6_and_42_ssc = core_wen & (and_777_rgt | and_779_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_781_rgt = and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1;
  assign and_783_rgt = and_dcpl_245 & and_dcpl_497;
  assign FpAdd_6U_10U_7_and_39_ssc = core_wen & (and_781_rgt | and_783_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_785_rgt = and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1;
  assign and_787_rgt = and_dcpl_245 & and_dcpl_501;
  assign FpAdd_6U_10U_7_and_40_ssc = core_wen & (and_785_rgt | and_787_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_789_rgt = and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1;
  assign and_791_rgt = and_dcpl_245 & and_dcpl_505;
  assign FpAdd_6U_10U_7_and_41_ssc = core_wen & (and_789_rgt | and_791_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign and_793_rgt = and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1;
  assign and_795_rgt = and_dcpl_245 & and_dcpl_509;
  assign FpAdd_6U_10U_7_and_42_ssc = core_wen & (and_793_rgt | and_795_rgt | and_dcpl_78)
      & mux_tmp_191;
  assign IsNaN_6U_10U_14_aelse_and_cse = core_wen & (~ and_dcpl_64) & mux_tmp_191;
  assign and_828_cse = or_181_cse & main_stage_v_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_cse = core_wen & (~ and_dcpl_64) &
      mux_tmp_192;
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_or_3_cse = and_dcpl_74 | and_dcpl_547;
  assign IsNaN_6U_10U_16_and_4_cse = core_wen & IsNaN_6U_10U_16_IsNaN_6U_10U_16_or_3_cse
      & mux_tmp_192;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_16_cse = core_wen & IsNaN_6U_10U_16_IsNaN_6U_10U_16_or_3_cse
      & mux_tmp_193;
  assign data_truncate_and_cse = core_wen & (~ and_dcpl_64) & mux_tmp_193;
  assign mux_194_nl = MUX_s_1_2_2(and_828_cse, mux_tmp_193, data_truncate_nor_dfs_4);
  assign and_2625_nl = data_truncate_nor_dfs_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt) & main_stage_v_4;
  assign mux_195_nl = MUX_s_1_2_2((and_2625_nl), (mux_194_nl), data_truncate_nor_dfs_3);
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_16_cse = core_wen & (~ and_dcpl_64)
      & (mux_195_nl);
  assign mux_196_nl = MUX_s_1_2_2(and_828_cse, mux_tmp_193, data_truncate_equal_tmp_4);
  assign and_2567_nl = data_truncate_equal_tmp_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt) & main_stage_v_4;
  assign mux_197_nl = MUX_s_1_2_2((and_2567_nl), (mux_196_nl), data_truncate_equal_tmp_3);
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_16_cse = core_wen & (~ and_dcpl_64)
      & (mux_197_nl);
  assign or_311_cse = IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_11_tmp | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  assign or_315_cse = data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_7_tmp;
  assign or_317_cse = (data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | IsNaN_6U_10U_16_land_4_lpi_1_dfm_3;
  assign nor_150_cse = ~((cfg_precision[0]) | (~ main_stage_v_1));
  assign and_2555_cse = or_tmp_302 & main_stage_v_4;
  assign nand_147_cse = ~((cfg_precision[1]) & or_181_cse);
  assign and_2550_cse = or_tmp_319 & main_stage_v_4;
  assign and_2545_cse = or_tmp_336 & main_stage_v_4;
  assign or_371_cse = data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_10_tmp;
  assign or_373_cse = data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_6_tmp;
  assign or_375_cse = data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_2_tmp;
  assign and_2537_cse = or_tmp_359 & main_stage_v_4;
  assign and_2532_cse = or_tmp_376 & main_stage_v_4;
  assign and_2527_cse = or_tmp_393 & main_stage_v_4;
  assign or_427_cse = IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_9_tmp | data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  assign or_429_cse = (data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | IsNaN_6U_10U_16_land_6_lpi_1_dfm_3;
  assign or_434_cse = (data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_2_lpi_1_dfm_3;
  assign and_2517_cse = or_tmp_419 & main_stage_v_4;
  assign and_2512_cse = or_tmp_441 & main_stage_v_4;
  assign or_476_cse = data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_8_tmp;
  assign and_2507_cse = data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign and_2503_cse = or_tmp_465 & main_stage_v_4;
  assign and_2498_cse = or_tmp_485 & main_stage_v_4;
  assign and_2491_cse = data_truncate_nor_tmp_4 & main_stage_v_3;
  assign and_2495_cse = main_stage_v_4 & data_truncate_nor_tmp_5;
  assign or_527_cse = and_2491_cse | m_row0_unequal_tmp_3 | (~ main_stage_v_2);
  assign or_521_cse = and_2491_cse | mux_tmp_364;
  assign and_2487_cse = or_tmp_513 & main_stage_v_4;
  assign or_548_cse = data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_14_tmp;
  assign and_2481_cse = or_tmp_532 & main_stage_v_4;
  assign or_567_cse = data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_13_tmp;
  assign and_2475_cse = or_tmp_551 & main_stage_v_4;
  assign and_2464_cse = or_tmp_579 & main_stage_v_4;
  assign IsNaN_6U_10U_16_and_cse = core_wen & (~((~ (cfg_precision[1])) | (~ main_stage_v_3)
      | and_dcpl_64));
  assign FpAdd_6U_10U_4_and_35_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_4_and_36_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_4_and_37_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_4_and_38_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_5_and_35_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_5_and_36_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_5_and_37_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_5_and_38_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_6_and_35_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_6_and_36_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_6_and_37_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_6_and_38_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_7_and_35_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_7_and_36_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_7_and_37_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1);
  assign FpAdd_6U_10U_7_and_38_ssc = core_wen & ((and_dcpl_245 & FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1
      & main_stage_v_2) | FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1);
  assign IsNaN_6U_10U_12_aelse_and_cse = core_wen & (~ or_dcpl_302);
  assign nand_nl = ~((~(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2619_nl = or_tmp_5 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_cse = MUX_s_1_2_2((and_2619_nl), (nand_nl), or_99_cse);
  assign and_932_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_645;
  assign and_935_rgt = and_dcpl_90 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_tmp);
  assign and_938_rgt = and_dcpl_99 & and_dcpl_94 & and_dcpl_651;
  assign and_941_rgt = and_dcpl_102 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_9_cse = core_wen & ((and_dcpl_74
      & and_dcpl_645) | and_dcpl_658) & mux_cse;
  assign nor_562_cse = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt);
  assign and_946_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_659;
  assign and_949_rgt = and_dcpl_120 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp);
  assign and_952_rgt = and_dcpl_129 & and_dcpl_124 & and_dcpl_665;
  assign and_955_rgt = and_dcpl_132 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
  assign or_14_nl = IsNaN_6U_10U_land_2_lpi_1_dfm | (~ or_dcpl_1);
  assign mux_3_nl = MUX_s_1_2_2(IsNaN_6U_10U_land_2_lpi_1_dfm, (or_14_nl), or_181_cse);
  assign mux_4_nl = MUX_s_1_2_2(IsNaN_6U_10U_land_2_lpi_1_dfm, (mux_3_nl), chn_data_in_rsci_bawt);
  assign or_15_nl = IsNaN_6U_10U_1_land_2_lpi_1_dfm | (mux_4_nl);
  assign mux_5_nl = MUX_s_1_2_2(IsNaN_6U_10U_land_2_lpi_1_dfm, and_72_cse, or_181_cse);
  assign mux_6_nl = MUX_s_1_2_2(IsNaN_6U_10U_land_2_lpi_1_dfm, (mux_5_nl), chn_data_in_rsci_bawt);
  assign mux_7_nl = MUX_s_1_2_2((mux_6_nl), nand_tmp_2, IsNaN_6U_10U_1_land_2_lpi_1_dfm);
  assign mux_8_nl = MUX_s_1_2_2((mux_7_nl), (or_15_nl), or_tmp_8);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_11_cse = core_wen & ((and_dcpl_74
      & and_dcpl_659) | and_dcpl_672) & (mux_8_nl);
  assign nand_3_nl = ~((~(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2618_nl = or_tmp_16 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_9_cse = MUX_s_1_2_2((and_2618_nl), (nand_3_nl), or_119_cse);
  assign and_960_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_673;
  assign and_963_rgt = and_dcpl_150 & and_dcpl_88 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp)
      & chn_data_in_rsci_bawt;
  assign and_966_rgt = and_dcpl_159 & and_dcpl_154 & and_dcpl_679;
  assign and_969_rgt = and_dcpl_162 & and_dcpl_88 & IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp
      & chn_data_in_rsci_bawt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse = core_wen & ((and_dcpl_74
      & and_dcpl_673) | and_dcpl_686) & mux_9_cse;
  assign nand_7_nl = ~((~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2616_nl = or_tmp_22 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_13_cse = MUX_s_1_2_2((and_2616_nl), (nand_7_nl), or_256_cse);
  assign and_974_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_687;
  assign and_977_rgt = and_dcpl_308 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign and_980_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_693;
  assign and_983_rgt = and_dcpl_90 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign and_985_rgt = and_dcpl_74 & and_dcpl_693;
  assign and_2462_nl = (~((~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35;
  assign nand_133_nl = ~(((~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp)
      & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_613_nl = (~ IsNaN_6U_10U_3_land_1_lpi_1_dfm) | IsNaN_6U_10U_2_land_1_lpi_1_dfm;
  assign mux_422_nl = MUX_s_1_2_2((nand_133_nl), (and_2462_nl), or_613_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse = core_wen & (~ or_dcpl_303)
      & (mux_422_nl);
  assign nand_11_nl = ~((~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2614_nl = or_tmp_25 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_16_cse = MUX_s_1_2_2((and_2614_nl), (nand_11_nl), or_237_cse);
  assign and_988_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_701;
  assign and_991_rgt = and_dcpl_282 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign and_994_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_707;
  assign and_997_rgt = and_dcpl_120 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign and_999_rgt = and_dcpl_74 & and_dcpl_707;
  assign and_2461_nl = (~((~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35;
  assign nand_132_nl = ~(((~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp)
      & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_615_nl = (~ IsNaN_6U_10U_3_land_2_lpi_1_dfm) | IsNaN_6U_10U_2_land_2_lpi_1_dfm;
  assign mux_423_nl = MUX_s_1_2_2((nand_132_nl), (and_2461_nl), or_615_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_2_cse = core_wen & (~ or_dcpl_303)
      & (mux_423_nl);
  assign and_1002_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_715;
  assign and_1005_rgt = and_dcpl_256 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign and_1008_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_721;
  assign and_1011_rgt = and_dcpl_150 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign and_1013_rgt = and_dcpl_74 & and_dcpl_721;
  assign and_2460_nl = (IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp | (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp))
      & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_424_nl = MUX_s_1_2_2(nand_tmp_61, (and_2460_nl), IsNaN_6U_10U_3_land_3_lpi_1_dfm);
  assign mux_425_nl = MUX_s_1_2_2((mux_424_nl), nand_tmp_61, IsNaN_6U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_4_cse = core_wen & (~ or_dcpl_303)
      & (~ (mux_425_nl));
  assign nand_23_nl = ~((~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2609_nl = or_tmp_33 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_27_cse = MUX_s_1_2_2((and_2609_nl), (nand_23_nl), or_209_cse);
  assign and_1016_rgt = and_dcpl_86 & and_dcpl_81 & and_dcpl_729;
  assign and_1019_rgt = and_dcpl_90 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
  assign and_1022_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_735;
  assign and_1025_rgt = and_dcpl_308 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_9_cse = core_wen & ((and_dcpl_74
      & and_dcpl_729) | and_dcpl_742) & mux_27_cse;
  assign nand_25_nl = ~((~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2608_nl = or_tmp_36 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_29_cse = MUX_s_1_2_2((and_2608_nl), (nand_25_nl), or_196_cse);
  assign and_1030_rgt = and_dcpl_117 & and_dcpl_112 & and_dcpl_743;
  assign and_1033_rgt = and_dcpl_120 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
  assign and_1036_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_749;
  assign and_1039_rgt = and_dcpl_282 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_10_cse = core_wen & ((and_dcpl_74
      & and_dcpl_743) | and_dcpl_756) & mux_29_cse;
  assign nand_27_nl = ~((~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2607_nl = or_tmp_39 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_31_cse = MUX_s_1_2_2((and_2607_nl), (nand_27_nl), or_183_cse);
  assign and_1044_rgt = and_dcpl_147 & and_dcpl_142 & and_dcpl_757;
  assign and_1047_rgt = and_dcpl_150 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign and_1050_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_763;
  assign and_1053_rgt = and_dcpl_256 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_11_cse = core_wen & ((and_dcpl_74
      & and_dcpl_757) | and_dcpl_770) & mux_31_cse;
  assign and_1058_rgt = and_dcpl_305 & and_dcpl_300 & and_dcpl_771;
  assign and_1061_rgt = and_dcpl_308 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign and_1064_rgt = and_dcpl_316 & and_dcpl_311 & and_dcpl_777;
  assign and_1067_rgt = and_dcpl_319 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign and_1069_rgt = and_dcpl_74 & and_dcpl_777;
  assign nand_33_nl = ~((~(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2605_nl = or_tmp_48 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_40_cse = MUX_s_1_2_2((and_2605_nl), (nand_33_nl), or_152_cse);
  assign and_1072_rgt = and_dcpl_279 & and_dcpl_274 & and_dcpl_785;
  assign and_1075_rgt = and_dcpl_282 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign and_1078_rgt = and_dcpl_290 & and_dcpl_285 & and_dcpl_791;
  assign and_1081_rgt = and_dcpl_293 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp);
  assign and_1083_rgt = and_dcpl_74 & and_dcpl_791;
  assign and_1086_rgt = and_dcpl_253 & and_dcpl_248 & and_dcpl_799;
  assign and_1089_rgt = and_dcpl_256 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign and_1092_rgt = and_dcpl_264 & and_dcpl_259 & and_dcpl_805;
  assign and_1095_rgt = and_dcpl_267 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign and_1097_rgt = and_dcpl_74 & and_dcpl_805;
  assign IsNaN_6U_10U_6_aelse_and_cse = core_wen & (~(or_dcpl_303 | (fsm_output[0])));
  assign FpAdd_6U_10U_3_b_int_mant_p1_and_cse = core_wen & (~ (fsm_output[0]));
  assign FpAdd_6U_10U_3_b_int_mant_p1_and_4_cse = FpAdd_6U_10U_3_b_int_mant_p1_and_cse
      & (~ or_dcpl_303);
  assign FpAdd_6U_10U_3_and_29_cse = core_wen & (and_1769_cse | and_1771_cse);
  assign or_617_nl = IsNaN_6U_10U_6_land_3_lpi_1_dfm | and_dcpl_52;
  assign and_125_nl = IsNaN_6U_10U_6_land_3_lpi_1_dfm & nand_tmp_2;
  assign mux_426_nl = MUX_s_1_2_2((and_125_nl), (or_617_nl), IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_12_cse = core_wen & (~ or_dcpl_303)
      & (mux_426_nl);
  assign FpAdd_6U_10U_3_and_32_cse = core_wen & (and_1801_cse | and_1803_cse);
  assign nand_63_nl = ~((~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2459_nl = IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_427_nl = MUX_s_1_2_2((and_2459_nl), (nand_63_nl), IsNaN_6U_10U_6_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_14_cse = core_wen & (~ or_dcpl_303)
      & (mux_427_nl);
  assign FpAdd_6U_10U_3_and_35_cse = core_wen & (and_1833_cse | and_1835_cse);
  assign mux_428_nl = MUX_s_1_2_2(and_tmp_1, or_tmp_45, IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_16_cse = core_wen & (~ or_dcpl_303)
      & (mux_428_nl);
  assign FpAdd_6U_10U_3_and_38_cse = core_wen & (and_1865_cse | and_1867_cse);
  assign FpAdd_6U_10U_2_and_29_cse = core_wen & (and_1895_cse | and_1897_cse);
  assign FpAdd_6U_10U_2_and_32_cse = core_wen & (and_1927_cse | and_1929_cse);
  assign FpAdd_6U_10U_2_and_35_cse = core_wen & (and_1959_cse | and_1961_cse);
  assign FpAdd_6U_10U_2_and_38_cse = core_wen & (and_1991_cse | and_1993_cse);
  assign FpAdd_6U_10U_1_and_29_cse = core_wen & (and_2021_cse | and_2023_cse);
  assign FpAdd_6U_10U_1_and_32_cse = core_wen & (and_2053_cse | and_2055_cse);
  assign FpAdd_6U_10U_1_and_35_cse = core_wen & (and_2085_cse | and_2087_cse);
  assign FpAdd_6U_10U_1_and_38_cse = core_wen & (and_2117_cse | and_2119_cse);
  assign FpAdd_6U_10U_and_29_cse = core_wen & (and_2147_cse | and_2149_cse);
  assign FpAdd_6U_10U_and_32_cse = core_wen & (and_2179_cse | and_2181_cse);
  assign FpAdd_6U_10U_and_35_cse = core_wen & (and_2211_cse | and_2213_cse);
  assign FpAdd_6U_10U_and_38_cse = core_wen & (and_2243_cse | and_2245_cse);
  assign or_623_cse = IsNaN_6U_10U_1_land_lpi_1_dfm | IsNaN_6U_10U_land_lpi_1_dfm_st;
  assign and_1268_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_975;
  assign and_1271_rgt = and_dcpl_985 & and_dcpl_88 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp);
  assign and_1280_rgt = and_dcpl_994 & and_dcpl_989 & and_dcpl_987;
  assign and_1283_rgt = and_dcpl_997 & and_dcpl_996;
  assign and_1285_rgt = or_dcpl_342 & or_181_cse;
  assign and_1288_rgt = or_dcpl_343 & or_181_cse;
  assign and_1291_rgt = (or_dcpl_1 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp) & or_181_cse;
  assign and_1294_rgt = or_dcpl_345 & or_181_cse;
  assign or_629_cse = IsNaN_6U_10U_7_land_lpi_1_dfm | IsNaN_6U_10U_6_land_lpi_1_dfm_st;
  assign and_1303_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1010;
  assign and_1306_rgt = and_dcpl_1020 & and_dcpl_1019;
  assign and_1314_rgt = and_dcpl_1028 & and_dcpl_1023 & and_dcpl_1007;
  assign and_1317_rgt = and_dcpl_1031 & and_dcpl_88 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_18_cse = core_wen & (and_dcpl_1033
      | and_dcpl_1034 | and_dcpl_1035) & mux_tmp_443;
  assign or_638_cse = IsNaN_6U_10U_5_land_lpi_1_dfm | IsNaN_6U_10U_4_land_lpi_1_dfm_st;
  assign and_1323_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_1036;
  assign and_1325_rgt = and_dcpl_985 & and_dcpl_88 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign and_1327_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1004;
  assign and_1329_rgt = and_dcpl_1020 & and_dcpl_88 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp);
  assign mux_447_nl = MUX_s_1_2_2(not_tmp_208, or_tmp_624, or_tmp_42);
  assign mux_448_nl = MUX_s_1_2_2(not_tmp_208, or_tmp_624, or_638_cse);
  assign mux_449_nl = MUX_s_1_2_2((mux_448_nl), (mux_447_nl), nor_57_cse);
  assign mux_450_nl = MUX_s_1_2_2(not_tmp_208, (mux_449_nl), chn_data_in_rsci_bawt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_18_cse = core_wen & (and_dcpl_1045
      | and_dcpl_78 | and_dcpl_1005) & (mux_450_nl);
  assign or_648_cse = IsNaN_6U_10U_3_land_lpi_1_dfm | IsNaN_6U_10U_2_land_lpi_1_dfm_st;
  assign and_1333_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1046;
  assign and_1335_rgt = and_dcpl_1020 & and_dcpl_1049;
  assign and_1337_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_1001;
  assign and_1339_rgt = and_dcpl_985 & and_dcpl_88 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_15_cse = core_wen & (and_dcpl_1055
      | and_dcpl_1002 | and_dcpl_1056) & mux_tmp_457;
  assign and_1342_rgt = and_dcpl_74 & and_dcpl_1046;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse = core_wen & (((~ mux_tmp_661)
      & or_181_cse) | and_dcpl_1059) & mux_tmp_460;
  assign and_1345_rgt = and_dcpl_74 & and_dcpl_987;
  assign mux_468_cse = MUX_s_1_2_2(main_stage_v_2, main_stage_v_1, or_181_cse);
  assign nor_592_nl = ~((~ main_stage_v_2) | (cfg_precision!=2'b00));
  assign mux_539_nl = MUX_s_1_2_2(main_stage_v_3, (nor_592_nl), or_181_cse);
  assign nor_593_nl = ~(nor_562_cse | (~ main_stage_v_2) | (cfg_precision!=2'b00));
  assign mux_540_nl = MUX_s_1_2_2((nor_593_nl), (mux_539_nl), data_truncate_equal_tmp_3);
  assign o_data_data_and_64_cse = core_wen & (~ and_dcpl_64) & (mux_540_nl);
  assign nor_445_nl = ~((~ main_stage_v_2) | (cfg_precision!=2'b01));
  assign mux_541_nl = MUX_s_1_2_2(main_stage_v_3, (nor_445_nl), or_181_cse);
  assign nor_446_nl = ~(nor_562_cse | (~ main_stage_v_2) | (cfg_precision!=2'b01));
  assign mux_542_nl = MUX_s_1_2_2((nor_446_nl), (mux_541_nl), data_truncate_nor_dfs_3);
  assign o_data_data_and_80_cse = core_wen & (~ and_dcpl_64) & (mux_542_nl);
  assign data_truncate_and_129_cse = (~ m_row0_unequal_tmp_3) & data_truncate_nor_tmp_mx0w0
      & (~ and_dcpl_64);
  assign data_truncate_and_130_cse = m_row0_unequal_tmp_3 & data_truncate_nor_tmp_mx0w0
      & (~ and_dcpl_64);
  assign data_truncate_data_truncate_nor_1_cse = ~((~(data_truncate_nor_dfs_mx0w0
      | data_truncate_equal_tmp_mx0w0)) | and_dcpl_64);
  assign data_truncate_and_124_cse = data_truncate_nor_dfs_mx0w0 & (~ and_dcpl_64);
  assign data_truncate_and_125_cse = data_truncate_equal_tmp_mx0w0 & (~ and_dcpl_64);
  assign nor_439_cse = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_12_land_1_lpi_1_dfm_4));
  assign or_796_cse = (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign or_840_nl = (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st;
  assign mux_571_nl = MUX_s_1_2_2(mux_tmp_570, or_tmp_823, or_840_nl);
  assign or_847_nl = (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st
      | or_tmp_828;
  assign nor_303_nl = ~(IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 | (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_5));
  assign mux_572_nl = MUX_s_1_2_2((or_847_nl), (mux_571_nl), nor_303_nl);
  assign FpAdd_6U_10U_2_o_expo_and_11_ssc = core_wen & (~ and_dcpl_64) & (~ (mux_572_nl));
  assign nor_387_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~((~((~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_3_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_3_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st)));
  assign nor_390_nl = ~((~((~(IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 | (~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_5)))
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_10_land_3_lpi_1_dfm_5))
      | (~ main_stage_v_3) | m_row0_unequal_tmp_4);
  assign mux_573_nl = MUX_s_1_2_2((nor_390_nl), (nor_387_nl), or_181_cse);
  assign FpAdd_6U_10U_2_o_expo_and_12_ssc = core_wen & (~ and_dcpl_64) & (mux_573_nl);
  assign or_856_nl = IsNaN_6U_10U_14_land_2_lpi_1_dfm_st | or_tmp_828;
  assign mux_574_nl = MUX_s_1_2_2(mux_tmp_570, or_tmp_823, IsNaN_6U_10U_14_land_2_lpi_1_dfm_st);
  assign or_855_nl = (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_2_lpi_1_dfm_5;
  assign mux_575_nl = MUX_s_1_2_2((mux_574_nl), (or_856_nl), or_855_nl);
  assign or_857_nl = (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_2_lpi_1_dfm_5
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_3) | m_row0_unequal_tmp_4;
  assign mux_576_nl = MUX_s_1_2_2((or_857_nl), (mux_575_nl), IsNaN_6U_10U_15_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_1_o_expo_and_11_ssc = core_wen & (~ and_dcpl_64) & (~ (mux_576_nl));
  assign nor_384_cse = ~(IsNaN_6U_10U_13_nor_1_itm_2 | IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2);
  assign nor_379_nl = ~((~ or_tmp_774) | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign nor_380_nl = ~((~(IsNaN_6U_10U_10_land_2_lpi_1_dfm_4 | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st))
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign nor_382_nl = ~((~(nor_384_cse | IsNaN_6U_10U_10_land_2_lpi_1_dfm_4 | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st))
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign or_861_nl = (cfg_precision!=2'b10) | IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3;
  assign mux_577_nl = MUX_s_1_2_2((nor_382_nl), (nor_380_nl), or_861_nl);
  assign mux_578_nl = MUX_s_1_2_2((mux_577_nl), (nor_379_nl), IsNaN_6U_10U_12_land_2_lpi_1_dfm_4);
  assign nor_385_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_11_land_2_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_13_land_2_lpi_1_dfm_3))) | IsNaN_6U_10U_14_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_2_lpi_1_dfm_5)));
  assign mux_579_nl = MUX_s_1_2_2((nor_385_nl), (mux_578_nl), or_181_cse);
  assign FpAdd_6U_10U_1_o_expo_and_12_ssc = core_wen & (~ and_dcpl_64) & (mux_579_nl);
  assign or_871_nl = IsNaN_6U_10U_14_land_1_lpi_1_dfm_st | or_tmp_828;
  assign mux_580_nl = MUX_s_1_2_2(mux_tmp_570, or_tmp_823, IsNaN_6U_10U_14_land_1_lpi_1_dfm_st);
  assign or_870_nl = (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_1_lpi_1_dfm_5;
  assign mux_581_nl = MUX_s_1_2_2((mux_580_nl), (or_871_nl), or_870_nl);
  assign or_872_nl = (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_1_lpi_1_dfm_5
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_3) | m_row0_unequal_tmp_4;
  assign mux_582_nl = MUX_s_1_2_2((or_872_nl), (mux_581_nl), IsNaN_6U_10U_15_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_o_expo_and_11_ssc = core_wen & (~ and_dcpl_64) & (~ (mux_582_nl));
  assign nor_374_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~((~((~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_1_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_1_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_1_lpi_1_dfm_st)));
  assign nor_377_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_9_land_1_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_5))) | IsNaN_6U_10U_14_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_1_lpi_1_dfm_5)));
  assign mux_583_nl = MUX_s_1_2_2((nor_377_nl), (nor_374_nl), or_181_cse);
  assign FpAdd_6U_10U_o_expo_and_12_ssc = core_wen & (~ and_dcpl_64) & (mux_583_nl);
  assign nor_370_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~(IsNaN_6U_10U_12_land_3_lpi_1_dfm_4
      | (~(IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 | or_tmp_738)))));
  assign nor_372_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_8_land_3_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_3))) | IsNaN_6U_10U_11_land_3_lpi_1_dfm_5)));
  assign mux_585_nl = MUX_s_1_2_2((nor_372_nl), (nor_370_nl), or_181_cse);
  assign FpAdd_6U_10U_2_o_expo_and_13_ssc = core_wen & (~ and_dcpl_64) & (mux_585_nl);
  assign nor_366_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~(IsNaN_6U_10U_12_land_2_lpi_1_dfm_4
      | (~(IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 | or_tmp_723)))));
  assign nor_368_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_8_land_2_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_3))) | IsNaN_6U_10U_11_land_2_lpi_1_dfm_5)));
  assign mux_587_nl = MUX_s_1_2_2((nor_368_nl), (nor_366_nl), or_181_cse);
  assign FpAdd_6U_10U_1_o_expo_and_13_ssc = core_wen & (~ and_dcpl_64) & (mux_587_nl);
  assign nor_364_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_5));
  assign mux_588_nl = MUX_s_1_2_2((nor_364_nl), nor_439_cse, or_181_cse);
  assign FpAdd_6U_10U_o_expo_and_13_ssc = core_wen & (~ and_dcpl_64) & (mux_588_nl);
  assign mux_589_nl = MUX_s_1_2_2(or_tmp_823, mux_tmp_570, IsNaN_6U_10U_8_land_3_lpi_1_dfm_4);
  assign nand_65_nl = ~(IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 & (~ or_tmp_828));
  assign mux_590_nl = MUX_s_1_2_2((nand_65_nl), (mux_589_nl), IsNaN_6U_10U_8_land_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_2_o_mant_and_8_cse = core_wen & (~ and_dcpl_64) & (~ (mux_590_nl));
  assign mux_591_nl = MUX_s_1_2_2(or_tmp_823, mux_tmp_570, IsNaN_6U_10U_8_land_2_lpi_1_dfm_4);
  assign nand_66_nl = ~(IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 & (~ or_tmp_828));
  assign mux_592_nl = MUX_s_1_2_2((nand_66_nl), (mux_591_nl), IsNaN_6U_10U_8_land_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_o_mant_and_8_cse = core_wen & (~ and_dcpl_64) & (~ (mux_592_nl));
  assign mux_593_nl = MUX_s_1_2_2(or_tmp_823, mux_tmp_570, IsNaN_6U_10U_8_land_1_lpi_1_dfm_4);
  assign nand_67_nl = ~(IsNaN_6U_10U_8_land_1_lpi_1_dfm_4 & (~ or_tmp_828));
  assign mux_594_nl = MUX_s_1_2_2((nand_67_nl), (mux_593_nl), IsNaN_6U_10U_8_land_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_o_mant_and_8_cse = core_wen & (~ and_dcpl_64) & (~ (mux_594_nl));
  assign or_917_nl = IsNaN_6U_10U_14_land_lpi_1_dfm_st | or_tmp_828;
  assign mux_595_nl = MUX_s_1_2_2(mux_tmp_570, or_tmp_823, IsNaN_6U_10U_14_land_lpi_1_dfm_st);
  assign or_916_nl = (~ IsNaN_6U_10U_15_land_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_lpi_1_dfm_5;
  assign mux_596_nl = MUX_s_1_2_2((mux_595_nl), (or_917_nl), or_916_nl);
  assign or_918_nl = (~ IsNaN_6U_10U_15_land_lpi_1_dfm_5) | IsNaN_6U_10U_14_land_lpi_1_dfm_5
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_3) | m_row0_unequal_tmp_4;
  assign mux_597_nl = MUX_s_1_2_2((or_918_nl), (mux_596_nl), IsNaN_6U_10U_15_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_3_o_expo_and_11_ssc = core_wen & (~ and_dcpl_64) & (~ (mux_597_nl));
  assign nor_355_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~((~((~ IsNaN_6U_10U_13_land_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_lpi_1_dfm_4 | IsNaN_6U_10U_14_land_lpi_1_dfm_st)));
  assign nor_358_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_11_land_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_13_land_lpi_1_dfm_5))) | IsNaN_6U_10U_14_land_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_lpi_1_dfm_5)));
  assign mux_598_nl = MUX_s_1_2_2((nor_358_nl), (nor_355_nl), or_181_cse);
  assign FpAdd_6U_10U_3_o_expo_and_12_ssc = core_wen & (~ and_dcpl_64) & (mux_598_nl);
  assign nor_351_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~(IsNaN_6U_10U_12_land_lpi_1_dfm_4
      | (~(IsNaN_6U_10U_8_land_lpi_1_dfm_4 | or_tmp_753)))));
  assign nor_353_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~((~(IsNaN_6U_10U_8_land_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_9_land_lpi_1_dfm_3))) | IsNaN_6U_10U_11_land_lpi_1_dfm_5)));
  assign mux_600_nl = MUX_s_1_2_2((nor_353_nl), (nor_351_nl), or_181_cse);
  assign FpAdd_6U_10U_3_o_expo_and_13_ssc = core_wen & (~ and_dcpl_64) & (mux_600_nl);
  assign mux_601_nl = MUX_s_1_2_2(or_tmp_823, mux_tmp_570, IsNaN_6U_10U_8_land_lpi_1_dfm_4);
  assign nand_68_nl = ~(IsNaN_6U_10U_8_land_lpi_1_dfm_4 & (~ or_tmp_828));
  assign mux_602_nl = MUX_s_1_2_2((nand_68_nl), (mux_601_nl), IsNaN_6U_10U_8_land_lpi_1_dfm_5);
  assign FpAdd_6U_10U_3_o_mant_and_8_cse = core_wen & (~ and_dcpl_64) & (~ (mux_602_nl));
  assign nand_5_nl = ~((~(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2617_nl = or_tmp_19 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_11_cse = MUX_s_1_2_2((and_2617_nl), (nand_5_nl), or_623_cse);
  assign and_1348_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_1061;
  assign and_1351_rgt = and_dcpl_985 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp);
  assign and_1354_rgt = and_dcpl_994 & and_dcpl_989 & and_dcpl_1067;
  assign and_1357_rgt = and_dcpl_997 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_18_cse = core_wen & ((and_dcpl_74
      & and_dcpl_1061) | and_dcpl_1074) & mux_11_cse;
  assign nand_19_nl = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2611_nl = or_tmp_30 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_24_cse = MUX_s_1_2_2((and_2611_nl), (nand_19_nl), or_648_cse);
  assign and_1362_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1075;
  assign and_1365_rgt = and_dcpl_1020 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  assign and_1368_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_1081;
  assign and_1371_rgt = and_dcpl_985 & and_dcpl_88 & chn_data_in_rsci_bawt & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign and_1373_rgt = and_dcpl_74 & and_dcpl_1081;
  assign and_2425_nl = (~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp | (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp)
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35;
  assign nand_123_nl = ~((IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp | (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp))
      & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_942_nl = (~ IsNaN_6U_10U_3_land_lpi_1_dfm) | IsNaN_6U_10U_2_land_lpi_1_dfm_st;
  assign mux_607_nl = MUX_s_1_2_2((nand_123_nl), (and_2425_nl), or_942_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse = core_wen & (~ or_dcpl_303)
      & (mux_607_nl);
  assign nand_29_nl = ~((~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2606_nl = or_tmp_42 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_33_cse = MUX_s_1_2_2((and_2606_nl), (nand_29_nl), or_638_cse);
  assign and_1376_rgt = and_dcpl_982 & and_dcpl_977 & and_dcpl_1089;
  assign and_1379_rgt = and_dcpl_985 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign and_1382_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1095;
  assign and_1385_rgt = and_dcpl_1020 & and_dcpl_88 & chn_data_in_rsci_bawt & (~
      IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_21_cse = core_wen & ((and_dcpl_74
      & and_dcpl_1089) | and_dcpl_1102) & mux_33_cse;
  assign nand_37_nl = ~((~(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign and_2603_nl = or_tmp_65 & chn_data_in_rsci_bawt & not_tmp_35;
  assign mux_46_cse = MUX_s_1_2_2((and_2603_nl), (nand_37_nl), or_629_cse);
  assign and_1390_rgt = and_dcpl_1017 & and_dcpl_1012 & and_dcpl_1103;
  assign and_1393_rgt = and_dcpl_1020 & and_dcpl_88 & chn_data_in_rsci_bawt & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign and_1396_rgt = and_dcpl_1028 & and_dcpl_1023 & and_dcpl_1109;
  assign and_1399_rgt = and_dcpl_1031 & and_dcpl_88 & chn_data_in_rsci_bawt & (~
      IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp);
  assign and_1401_rgt = and_dcpl_74 & and_dcpl_1109;
  assign nand_71_nl = ~((~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2424_nl = IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_608_nl = MUX_s_1_2_2((and_2424_nl), (nand_71_nl), IsNaN_6U_10U_6_land_lpi_1_dfm_st);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_22_cse = core_wen & (~ or_dcpl_303)
      & (mux_608_nl);
  assign FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse = and_dcpl_1119 | and_dcpl_1122;
  assign mux_629_nl = MUX_s_1_2_2(IsNaN_6U_10U_8_land_2_lpi_1_dfm_st, IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp,
      nor_57_cse);
  assign and_2423_nl = main_stage_v_1 & (~ (mux_629_nl));
  assign nor_349_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3);
  assign mux_630_nl = MUX_s_1_2_2((nor_349_nl), (and_2423_nl), or_181_cse);
  assign IsNaN_6U_10U_9_and_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & (mux_630_nl);
  assign mux_631_nl = MUX_s_1_2_2(IsNaN_6U_10U_8_land_3_lpi_1_dfm_st, IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp,
      nor_57_cse);
  assign and_2422_nl = main_stage_v_1 & (~ (mux_631_nl));
  assign nor_348_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3);
  assign mux_632_nl = MUX_s_1_2_2((nor_348_nl), (and_2422_nl), or_181_cse);
  assign IsNaN_6U_10U_9_and_7_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & (mux_632_nl);
  assign mux_633_nl = MUX_s_1_2_2(IsNaN_6U_10U_8_land_lpi_1_dfm_st, IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp,
      nor_57_cse);
  assign and_2421_nl = main_stage_v_1 & (~ (mux_633_nl));
  assign nor_347_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_8_land_lpi_1_dfm_st_3);
  assign mux_634_nl = MUX_s_1_2_2((nor_347_nl), (and_2421_nl), or_181_cse);
  assign IsNaN_6U_10U_9_and_9_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & (mux_634_nl);
  assign mux_635_nl = MUX_s_1_2_2(or_tmp_976, IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp,
      or_181_cse);
  assign nor_346_nl = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ or_tmp_976));
  assign mux_636_nl = MUX_s_1_2_2((nor_346_nl), or_tmp_977, IsNaN_6U_10U_12_land_2_lpi_1_dfm_st);
  assign mux_637_nl = MUX_s_1_2_2((mux_636_nl), (mux_635_nl), nor_57_cse);
  assign mux_638_nl = MUX_s_1_2_2(or_tmp_977, (mux_637_nl), main_stage_v_1);
  assign IsNaN_6U_10U_13_and_cse = core_wen & IsNaN_6U_10U_6_aelse_IsNaN_6U_10U_6_aelse_or_7_cse
      & (~ (mux_638_nl));
  assign IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse = or_dcpl_366 & (~ and_dcpl_64);
  assign IntShiftRight_18U_2U_16U_mbits_fixed_and_cse = core_wen & ((~(or_dcpl_366
      | and_dcpl_64)) | IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse) & mux_468_cse;
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_80_cse = core_wen & (((cfg_precision==2'b01)
      & or_181_cse) | and_dcpl_1126) & mux_468_cse;
  assign IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse = or_dcpl_367 & (~ and_dcpl_64);
  assign IntShiftRight_18U_2U_8U_mbits_fixed_and_cse = core_wen & ((~(or_dcpl_367
      | and_dcpl_64)) | IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse) & mux_468_cse;
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_144_cse = core_wen & (((cfg_precision==2'b00)
      & or_181_cse) | and_dcpl_1129) & mux_468_cse;
  assign FpAdd_6U_10U_o_sign_or_1_rgt = (or_181_cse & and_dcpl_1131) | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp)
      & FpAdd_6U_10U_o_sign_1_lpi_1_dfm_3_mx0c2);
  assign FpAdd_6U_10U_1_o_sign_or_1_rgt = (or_181_cse & and_dcpl_1136) | ((~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp)
      & FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_3_mx0c2);
  assign nor_345_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp | or_tmp_966);
  assign nand_118_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp & (~ or_tmp_966));
  assign mux_645_nl = MUX_s_1_2_2((nand_118_nl), (nor_345_nl), IsNaN_6U_10U_8_land_2_lpi_1_dfm_st);
  assign IsNaN_6U_10U_9_and_11_cse = FpAdd_6U_10U_3_b_int_mant_p1_and_cse & (~ or_dcpl_302)
      & (mux_645_nl);
  assign m_row1_if_d2_or_1_rgt = (or_181_cse & and_dcpl_1141) | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp)
      & FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_3_mx0c2);
  assign nor_344_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp | or_tmp_966);
  assign nand_117_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp & (~ or_tmp_966));
  assign mux_646_nl = MUX_s_1_2_2((nand_117_nl), (nor_344_nl), IsNaN_6U_10U_8_land_3_lpi_1_dfm_st);
  assign IsNaN_6U_10U_9_and_13_cse = FpAdd_6U_10U_3_b_int_mant_p1_and_cse & (~ or_dcpl_302)
      & (mux_646_nl);
  assign FpAdd_6U_10U_1_o_sign_or_4_rgt = (or_181_cse & and_dcpl_1146) | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp)
      & FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_3_mx0c2);
  assign nor_343_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp | or_tmp_966);
  assign nand_116_nl = ~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp & (~ or_tmp_966));
  assign mux_647_nl = MUX_s_1_2_2((nand_116_nl), (nor_343_nl), IsNaN_6U_10U_8_land_lpi_1_dfm_st);
  assign IsNaN_6U_10U_9_and_15_cse = FpAdd_6U_10U_3_b_int_mant_p1_and_cse & (~ or_dcpl_302)
      & (mux_647_nl);
  assign and_1439_m1c = or_181_cse & and_dcpl_1153;
  assign FpAdd_6U_10U_o_sign_or_11_rgt = (or_181_cse & and_dcpl_1151) | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp)
      & and_1439_m1c);
  assign and_1440_rgt = or_181_cse & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign and_1442_rgt = or_181_cse & and_dcpl_1156;
  assign and_1444_rgt = or_181_cse & and_dcpl_1158;
  assign and_1449_m1c = or_181_cse & and_dcpl_1163;
  assign m_row1_if_d2_or_11_rgt = (or_181_cse & and_dcpl_1161) | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp)
      & and_1449_m1c);
  assign and_1454_m1c = or_181_cse & and_dcpl_1168;
  assign FpAdd_6U_10U_1_o_sign_or_17_rgt = (or_181_cse & and_dcpl_1166) | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp)
      & and_1454_m1c);
  assign and_1459_m1c = or_181_cse & and_dcpl_1173;
  assign FpAdd_6U_10U_o_sign_or_8_rgt = (or_181_cse & and_dcpl_1171) | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp)
      & and_1459_m1c);
  assign and_1460_rgt = or_181_cse & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign and_1462_rgt = or_181_cse & and_dcpl_1176;
  assign and_1464_rgt = or_181_cse & and_dcpl_1178;
  assign nor_342_nl = ~(IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp | or_tmp_966);
  assign nand_115_nl = ~(IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp & (~ or_tmp_966));
  assign mux_648_nl = MUX_s_1_2_2((nand_115_nl), (nor_342_nl), IsNaN_6U_10U_12_land_2_lpi_1_dfm_st);
  assign IsNaN_6U_10U_13_and_3_cse = FpAdd_6U_10U_3_b_int_mant_p1_and_cse & (~ or_dcpl_302)
      & (mux_648_nl);
  assign and_1469_m1c = or_181_cse & and_dcpl_1183;
  assign m_row1_if_d2_or_8_rgt = (or_181_cse & and_dcpl_1181) | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp)
      & and_1469_m1c);
  assign and_1474_m1c = or_181_cse & and_dcpl_1188;
  assign FpAdd_6U_10U_1_o_sign_or_14_rgt = (or_181_cse & and_dcpl_1186) | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp)
      & and_1474_m1c);
  assign FpAdd_6U_10U_1_o_sign_or_9_rgt = (or_181_cse & and_dcpl_1191) | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp)
      & FpAdd_6U_10U_3_o_sign_lpi_1_dfm_3_mx0c2);
  assign m_row1_if_d2_or_3_rgt = (or_181_cse & and_dcpl_1196) | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp)
      & FpAdd_6U_10U_2_o_sign_lpi_1_dfm_3_mx0c2);
  assign FpAdd_6U_10U_1_o_sign_or_6_rgt = (or_181_cse & and_dcpl_1201) | ((~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp)
      & FpAdd_6U_10U_1_o_sign_lpi_1_dfm_3_mx0c2);
  assign FpAdd_6U_10U_o_sign_or_3_rgt = (or_181_cse & and_dcpl_1206) | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp)
      & FpAdd_6U_10U_o_sign_lpi_1_dfm_3_mx0c2);
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_cse = core_wen & (~(or_dcpl_368
      | (~ (cfg_precision[0])) | and_dcpl_64));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_cse = core_wen & (~(or_dcpl_368
      | (cfg_precision[0]) | and_dcpl_64));
  assign IntSubExt_16U_16U_17U_2_o_and_cse = core_wen & (~(and_dcpl_88 | and_dcpl_64
      | (~ chn_data_in_rsci_bawt) | (fsm_output[0])));
  assign and_337_nl = and_dcpl_52 & (fsm_output[1]);
  assign m_row3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln477_assert_iExpoWidth_le_oExpoWidth_7_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_337_nl);
  assign and_339_nl = or_dcpl_1 & or_181_cse & chn_data_in_rsci_bawt & (fsm_output[1]);
  assign o_col3_4_NV_NVDLA_CSC_pra_cell_core_nvdla_int_h_ln274_assert_oWidth_gt_mWidth_5_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_339_nl);
  assign or_1110_nl = (or_181_cse & (cfg_precision[1]) & chn_data_in_rsci_bawt &
      (fsm_output[1])) | ((cfg_precision[1]) & chn_data_out_rsci_bawt & and_dcpl_57);
  assign data_truncate_16_NV_NVDLA_CSC_pra_cell_core_nvdla_float_h_ln630_assert_iExpoWidth_gt_oExpoWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, or_1110_nl);
  assign IsZero_5U_10U_1_aelse_not_18_nl = ~ IsZero_5U_10U_1_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[137:128]), (IsZero_5U_10U_1_aelse_not_18_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_33_nl = MUX_v_10_2_2(m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_33_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl = MUX_v_10_2_2(10'b0000000000,
      (chn_data_in_rsci_d_mxwt[9:0]), IsZero_5U_10U_aelse_not_19);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl = MUX_v_10_2_2(m_row0_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w4 =
      MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl), 10'b1111111111, IsInf_5U_10U_land_1_lpi_1_dfm);
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp = m_row0_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsZero_5U_10U_1_aelse_not_16_nl = ~ IsZero_5U_10U_1_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[153:144]), (IsZero_5U_10U_1_aelse_not_16_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_37_nl = MUX_v_10_2_2(m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_3_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_37_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[25:16]), IsZero_5U_10U_aelse_not_17);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_24_nl = MUX_v_10_2_2(m_row0_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_2_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_24_nl), 10'b1111111111,
      IsInf_5U_10U_land_2_lpi_1_dfm);
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp = m_row0_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsZero_5U_10U_1_aelse_not_14_nl = ~ IsZero_5U_10U_1_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_6_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[169:160]), (IsZero_5U_10U_1_aelse_not_14_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_31_nl = MUX_v_10_2_2(m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_31_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[41:32]), IsZero_5U_10U_aelse_not_15);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_25_nl = MUX_v_10_2_2(m_row0_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_25_nl), 10'b1111111111,
      IsInf_5U_10U_land_3_lpi_1_dfm);
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp = m_row0_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp = m_row0_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp = m_row0_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp = m_row0_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp = m_row2_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp = m_row2_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp = m_row2_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2==4'b1111);
  assign IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2==4'b1111);
  assign IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2==4'b1111);
  assign m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[127]) ^ (chn_data_in_rsci_d_mxwt[255]);
  assign nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign nl_FpAdd_6U_10U_3_is_a_greater_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_3_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_3_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_3_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0}) != ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2})))) | (readslicef_7_1_6((FpAdd_6U_10U_3_is_a_greater_acc_3_nl)));
  assign IsZero_5U_10U_2_aelse_not_14_nl = ~ IsZero_5U_10U_2_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_6_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[105:96]), (IsZero_5U_10U_2_aelse_not_14_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_31_nl = MUX_v_10_2_2(m_row1_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_31_nl), 10'b1111111111,
      IsInf_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_6_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[233:224]), IsZero_5U_10U_7_aelse_not_15);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_25_nl = MUX_v_10_2_2(m_row3_3_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_4_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_25_nl), 10'b1111111111,
      IsInf_5U_10U_7_land_3_lpi_1_dfm);
  assign IsZero_5U_10U_2_aelse_not_22_nl = ~ IsZero_5U_10U_2_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_8_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[109:106]), (IsZero_5U_10U_2_aelse_not_22_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_cse
      , IsDenorm_5U_10U_2_land_3_lpi_1_dfm , IsInf_5U_10U_2_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl),
      4'b1111, IsNaN_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_8_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[237:234]), IsZero_5U_10U_7_aelse_not_15);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_2_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_2_cse
      , IsDenorm_5U_10U_7_land_3_lpi_1_dfm , IsInf_5U_10U_7_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_2_nl),
      4'b1111, IsNaN_5U_10U_7_land_3_lpi_1_dfm);
  assign m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[111]) ^ (chn_data_in_rsci_d_mxwt[239]);
  assign nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign nl_FpAdd_6U_10U_3_is_a_greater_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_3_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_3_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_2_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) != ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2})))) | (readslicef_7_1_6((FpAdd_6U_10U_3_is_a_greater_acc_2_nl)));
  assign IsZero_5U_10U_2_aelse_not_16_nl = ~ IsZero_5U_10U_2_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[89:80]), (IsZero_5U_10U_2_aelse_not_16_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_35_nl = MUX_v_10_2_2(m_row1_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_3_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_35_nl), 10'b1111111111,
      IsInf_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[217:208]), IsZero_5U_10U_7_aelse_not_17);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_24_nl = MUX_v_10_2_2(m_row3_2_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_3_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_2_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_24_nl), 10'b1111111111,
      IsInf_5U_10U_7_land_2_lpi_1_dfm);
  assign IsZero_5U_10U_2_aelse_not_24_nl = ~ IsZero_5U_10U_2_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_5_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[93:90]), (IsZero_5U_10U_2_aelse_not_24_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_cse
      , IsDenorm_5U_10U_2_land_2_lpi_1_dfm , IsInf_5U_10U_2_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl),
      4'b1111, IsNaN_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_5_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[221:218]), IsZero_5U_10U_7_aelse_not_17);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_1_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_1_cse
      , IsDenorm_5U_10U_7_land_2_lpi_1_dfm , IsInf_5U_10U_7_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_1_nl),
      4'b1111, IsNaN_5U_10U_7_land_2_lpi_1_dfm);
  assign m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[95]) ^ (chn_data_in_rsci_d_mxwt[223]);
  assign nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign nl_FpAdd_6U_10U_3_is_a_greater_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_3_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_3_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_1_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) != ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2})))) | (readslicef_7_1_6((FpAdd_6U_10U_3_is_a_greater_acc_1_nl)));
  assign IsZero_5U_10U_2_aelse_not_18_nl = ~ IsZero_5U_10U_2_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[73:64]), (IsZero_5U_10U_2_aelse_not_18_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_37_nl = MUX_v_10_2_2(m_row1_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_37_nl), 10'b1111111111,
      IsInf_5U_10U_2_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[201:192]), IsZero_5U_10U_7_aelse_not_19);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_26_nl = MUX_v_10_2_2(m_row3_1_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_26_nl), 10'b1111111111,
      IsInf_5U_10U_7_land_1_lpi_1_dfm);
  assign IsZero_5U_10U_2_aelse_not_26_nl = ~ IsZero_5U_10U_2_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_2_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[77:74]), (IsZero_5U_10U_2_aelse_not_26_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_cse
      , IsDenorm_5U_10U_2_land_1_lpi_1_dfm , IsInf_5U_10U_2_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl),
      4'b1111, IsNaN_5U_10U_2_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_2_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[205:202]), IsZero_5U_10U_7_aelse_not_19);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_cse
      , IsDenorm_5U_10U_7_land_1_lpi_1_dfm , IsInf_5U_10U_7_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_nl),
      4'b1111, IsNaN_5U_10U_7_land_1_lpi_1_dfm);
  assign m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[79]) ^ (chn_data_in_rsci_d_mxwt[207]);
  assign nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl[10:0];
  assign nl_FpAdd_6U_10U_3_is_a_greater_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_3_is_a_greater_acc_nl = nl_FpAdd_6U_10U_3_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_3_is_a_greater_oif_aelse_acc_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) != ({FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2})))) | (readslicef_7_1_6((FpAdd_6U_10U_3_is_a_greater_acc_nl)));
  assign m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[191]) ^ (chn_data_in_rsci_d_mxwt[127]);
  assign nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign nl_FpAdd_6U_10U_2_is_a_greater_acc_3_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_2_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_2_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_3_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_2_is_a_greater_acc_3_nl)));
  assign IsZero_5U_10U_1_aelse_not_22_nl = ~ IsZero_5U_10U_1_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_8_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[173:170]), (IsZero_5U_10U_1_aelse_not_22_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_8_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse
      , IsDenorm_5U_10U_1_land_3_lpi_1_dfm , IsInf_5U_10U_1_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_8_nl),
      4'b1111, IsNaN_5U_10U_1_land_3_lpi_1_dfm);
  assign m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[175]) ^ (chn_data_in_rsci_d_mxwt[111]);
  assign nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , m_row2_if_d1_mux_7_cse})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign nl_FpAdd_6U_10U_2_is_a_greater_acc_2_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_2_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_2_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_2_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_2_is_a_greater_acc_2_nl)));
  assign IsZero_5U_10U_1_aelse_not_24_nl = ~ IsZero_5U_10U_1_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_5_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[157:154]), (IsZero_5U_10U_1_aelse_not_24_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_6_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse
      , IsDenorm_5U_10U_1_land_2_lpi_1_dfm , IsInf_5U_10U_1_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_6_nl),
      4'b1111, IsNaN_5U_10U_1_land_2_lpi_1_dfm);
  assign m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[159]) ^ (chn_data_in_rsci_d_mxwt[95]);
  assign nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , m_row2_if_d1_mux_4_cse})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign nl_FpAdd_6U_10U_2_is_a_greater_acc_1_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_2_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_2_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_1_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_2_is_a_greater_acc_1_nl)));
  assign IsZero_5U_10U_1_aelse_not_26_nl = ~ IsZero_5U_10U_1_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_2_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[141:138]), (IsZero_5U_10U_1_aelse_not_26_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_4_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse
      , IsDenorm_5U_10U_1_land_1_lpi_1_dfm , IsInf_5U_10U_1_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_4_nl),
      4'b1111, IsNaN_5U_10U_1_land_1_lpi_1_dfm);
  assign m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[143]) ^ (chn_data_in_rsci_d_mxwt[79]);
  assign nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl = ({1'b1 , m_row2_if_d1_mux_1_cse})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0)
      + 11'b1;
  assign FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl[10:0];
  assign nl_FpAdd_6U_10U_2_is_a_greater_acc_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)}) + 7'b1;
  assign FpAdd_6U_10U_2_is_a_greater_acc_nl = nl_FpAdd_6U_10U_2_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_2_is_a_greater_oif_aelse_acc_nl)))
      | (({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_2_is_a_greater_acc_nl)));
  assign m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~((chn_data_in_rsci_d_mxwt[127]) ^ (chn_data_in_rsci_d_mxwt[191]));
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1)
      + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0)})
      + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0})
      != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_3_nl)));
  assign IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp = m_row2_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~((chn_data_in_rsci_d_mxwt[111]) ^ (chn_data_in_rsci_d_mxwt[175]));
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_7_cse) + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0)})
      + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0})
      != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_2_nl)));
  assign IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp = m_row2_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~((chn_data_in_rsci_d_mxwt[95]) ^ (chn_data_in_rsci_d_mxwt[159]));
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_4_cse) + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0)})
      + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0})
      != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_1_nl)));
  assign IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp = m_row2_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~((chn_data_in_rsci_d_mxwt[79]) ^ (chn_data_in_rsci_d_mxwt[143]));
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_1_cse) + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl[10:0];
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_nl = ({1'b1 , (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0)})
      + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0})
      != ({(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]) , FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0})))) | (readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_nl)));
  assign m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[63]) ^ (chn_data_in_rsci_d_mxwt[191]);
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1)
      + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign nl_FpAdd_6U_10U_is_a_greater_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2})
      != ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0}))))
      | (readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_3_nl)));
  assign IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2==4'b1111);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl =
      MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[45:42]), IsZero_5U_10U_aelse_not_15);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse
      , IsDenorm_5U_10U_land_3_lpi_1_dfm , IsInf_5U_10U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl),
      4'b1111, IsNaN_5U_10U_land_3_lpi_1_dfm);
  assign m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[47]) ^ (chn_data_in_rsci_d_mxwt[175]);
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_7_cse) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign nl_FpAdd_6U_10U_is_a_greater_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2})
      != ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0}))))
      | (readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_2_nl)));
  assign IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2==4'b1111);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl =
      MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[29:26]), IsZero_5U_10U_aelse_not_17);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse
      , IsDenorm_5U_10U_land_2_lpi_1_dfm , IsInf_5U_10U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl),
      4'b1111, IsNaN_5U_10U_land_2_lpi_1_dfm);
  assign m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[31]) ^ (chn_data_in_rsci_d_mxwt[159]);
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_4_cse) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign nl_FpAdd_6U_10U_is_a_greater_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2})
      != ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0}))))
      | (readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_1_nl)));
  assign IsNaN_6U_10U_IsNaN_6U_10U_and_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2==4'b1111);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl =
      MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[13:10]), IsZero_5U_10U_aelse_not_19);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse
      , IsDenorm_5U_10U_land_1_lpi_1_dfm , IsInf_5U_10U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl),
      4'b1111, IsNaN_5U_10U_land_1_lpi_1_dfm);
  assign m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0
      = (chn_data_in_rsci_d_mxwt[15]) ^ (chn_data_in_rsci_d_mxwt[143]);
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0})
      + conv_u2u_10_11(~ m_row2_if_d1_mux_1_cse) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl[10:0];
  assign nl_FpAdd_6U_10U_is_a_greater_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4
      , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}) + conv_u2u_6_7({(~
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_nl = nl_FpAdd_6U_10U_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp = (~((readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl)))
      | (({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2})
      != ({FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4 , FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0}))))
      | (readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_nl)));
  assign o_col0_1_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col0_2_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col0_3_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col0_4_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col1_1_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col1_2_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col1_3_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col1_4_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2});
  assign o_col2_1_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2});
  assign o_col2_2_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2});
  assign o_col2_3_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2});
  assign o_col2_4_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2});
  assign o_col3_1_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2});
  assign o_col3_2_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2});
  assign o_col3_3_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2});
  assign o_col3_4_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp = ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2})
      == ({reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2});
  assign nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_4_o_expo_1_lpi_2)}) + 7'b10001;
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_4_o_expo_1_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_5_o_expo_1_lpi_2)}) + 7'b10001;
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_5_o_expo_1_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_6_o_expo_1_lpi_2)}) + 7'b10001;
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_6_o_expo_1_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_7_o_expo_1_lpi_2)}) + 7'b10001;
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_7_o_expo_1_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_4_o_expo_2_lpi_2)}) + 7'b10001;
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_4_o_expo_2_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_5_o_expo_2_lpi_2)}) + 7'b10001;
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_5_o_expo_2_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_6_o_expo_2_lpi_2)}) + 7'b10001;
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_6_o_expo_2_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_7_o_expo_2_lpi_2)}) + 7'b10001;
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_7_o_expo_2_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_4_o_expo_3_lpi_2)}) + 7'b10001;
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 = readslicef_7_1_6((data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_4_o_expo_3_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_5_o_expo_3_lpi_2)}) + 7'b10001;
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_5_o_expo_3_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_6_o_expo_3_lpi_2)}) + 7'b10001;
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_6_o_expo_3_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_7_o_expo_3_lpi_2)}) + 7'b10001;
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_7_o_expo_3_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_4_o_expo_lpi_2)}) + 7'b10001;
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_4_o_expo_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_5_o_expo_lpi_2)}) + 7'b10001;
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_5_o_expo_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_6_o_expo_lpi_2)}) + 7'b10001;
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_6_o_expo_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_6U_10U_7_o_expo_lpi_2)}) + 7'b10001;
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl = nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl[6:0];
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1 =
      readslicef_7_1_6((data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_5_6(FpAdd_6U_10U_7_o_expo_lpi_2[5:1])
      + 6'b111101;
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl = nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl[5:0];
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1 = readslicef_6_1_5((data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_7_o_expo_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_nor_15_tmp = ~((FpAdd_6U_10U_7_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_tmp = ~((FpAdd_6U_10U_7_o_expo_lpi_1_dfm_8_mx0w0==6'b111111));
  assign nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_6_o_expo_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_14_tmp = ~((~((FpAdd_6U_10U_6_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_6_o_expo_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_5_o_expo_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_13_tmp = ~((~((FpAdd_6U_10U_5_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_5_o_expo_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_4_o_expo_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_nor_12_tmp = ~((FpAdd_6U_10U_4_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_tmp = ~((FpAdd_6U_10U_4_o_expo_lpi_1_dfm_8_mx0w0==6'b111111));
  assign nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_11_tmp = ~((~((FpAdd_6U_10U_7_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_10_tmp = ~((~((FpAdd_6U_10U_6_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_9_tmp = ~((~((FpAdd_6U_10U_5_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_8_tmp = ~((~((FpAdd_6U_10U_4_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_7_tmp = ~((~((FpAdd_6U_10U_7_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_6_tmp = ~((~((FpAdd_6U_10U_6_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_5_tmp = ~((~((FpAdd_6U_10U_5_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_4_tmp = ~((~((FpAdd_6U_10U_4_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_3_tmp = ~((~((FpAdd_6U_10U_7_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_2_tmp = ~((~((FpAdd_6U_10U_6_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_1_tmp = ~((~((FpAdd_6U_10U_5_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = conv_u2s_6_7(FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_8_mx0w0)
      + 7'b1010001;
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl = nl_data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl[6:0];
  assign data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 = readslicef_7_1_6((data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_nl));
  assign IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_tmp = ~((~((FpAdd_6U_10U_4_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_8_mx0w0!=6'b111111));
  assign m_row0_m_row0_nor_15_m1c = ~(IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl = (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_7_else_carry_3_sva);
  assign o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl = nl_o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl[9:0];
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_10_nl = MUX_v_10_2_2((o_col3_3_FpMantRNE_23U_11U_7_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0);
  assign m_row0_and_49_nl = (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_5) & m_row0_m_row0_nor_15_m1c;
  assign m_row0_and_50_nl = IsNaN_6U_10U_15_land_3_lpi_1_dfm_5 & m_row0_m_row0_nor_15_m1c;
  assign FpAdd_6U_10U_7_o_mant_3_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_10_nl),
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_7, FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_7_o_mant_3_lpi_2,
      {(m_row0_and_49_nl) , (m_row0_and_50_nl) , m_row0_asn_184 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_14_m1c = ~(IsNaN_6U_10U_14_land_2_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl = (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_7_else_carry_2_sva);
  assign o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl = nl_o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl[9:0];
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_9_nl = MUX_v_10_2_2((o_col3_2_FpMantRNE_23U_11U_7_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0);
  assign m_row0_and_51_nl = (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_5) & m_row0_m_row0_nor_14_m1c;
  assign m_row0_and_52_nl = IsNaN_6U_10U_15_land_2_lpi_1_dfm_5 & m_row0_m_row0_nor_14_m1c;
  assign FpAdd_6U_10U_7_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_9_nl),
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_7, FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_7_o_mant_2_lpi_2,
      {(m_row0_and_51_nl) , (m_row0_and_52_nl) , m_row0_asn_186 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_13_m1c = ~(IsNaN_6U_10U_14_land_1_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl = (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_7_else_carry_1_sva);
  assign o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl = nl_o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl[9:0];
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_8_nl = MUX_v_10_2_2((o_col3_1_FpMantRNE_23U_11U_7_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0);
  assign m_row0_and_53_nl = (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_5) & m_row0_m_row0_nor_13_m1c;
  assign m_row0_and_54_nl = IsNaN_6U_10U_15_land_1_lpi_1_dfm_5 & m_row0_m_row0_nor_13_m1c;
  assign FpAdd_6U_10U_7_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_8_nl),
      FpAdd_6U_10U_o_mant_lpi_1_dfm_7, FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_7_o_mant_1_lpi_2,
      {(m_row0_and_53_nl) , (m_row0_and_54_nl) , m_row0_asn_188 , m_row0_unequal_tmp_4});
  assign nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl = FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_2
      + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl = nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_31_nl = (~(FpAdd_6U_10U_7_and_2_tmp | FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_19_nl = FpAdd_6U_10U_7_and_2_tmp & (~ FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_32_nl = FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_9_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_21_nl = IsNaN_6U_10U_15_land_3_lpi_1_dfm_5 & (~ IsNaN_6U_10U_14_land_3_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_2,
      (o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_7_o_expo_3_lpi_2,
      {(FpAdd_6U_10U_7_and_31_nl) , (FpAdd_6U_10U_7_and_19_nl) , (FpAdd_6U_10U_7_and_32_nl)
      , (FpAdd_6U_10U_7_and_21_nl) , m_row0_asn_184 , m_row0_unequal_tmp_4});
  assign nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl = FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_2
      + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl = nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_29_nl = (~(FpAdd_6U_10U_7_and_1_tmp | FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_13_nl = FpAdd_6U_10U_7_and_1_tmp & (~ FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_30_nl = FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_7_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_15_nl = IsNaN_6U_10U_15_land_2_lpi_1_dfm_5 & (~ IsNaN_6U_10U_14_land_2_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_2,
      (o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_7_o_expo_2_lpi_2,
      {(FpAdd_6U_10U_7_and_29_nl) , (FpAdd_6U_10U_7_and_13_nl) , (FpAdd_6U_10U_7_and_30_nl)
      , (FpAdd_6U_10U_7_and_15_nl) , m_row0_asn_186 , m_row0_unequal_tmp_4});
  assign nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl = FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_2
      + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl = nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_nl = (~(FpAdd_6U_10U_7_and_tmp | FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_6_nl = FpAdd_6U_10U_7_and_tmp & (~ FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_28_nl = FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_5_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_9_nl = IsNaN_6U_10U_15_land_1_lpi_1_dfm_5 & (~ IsNaN_6U_10U_14_land_1_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_2,
      (o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_7_o_expo_1_lpi_2,
      {(FpAdd_6U_10U_7_and_nl) , (FpAdd_6U_10U_7_and_6_nl) , (FpAdd_6U_10U_7_and_28_nl)
      , (FpAdd_6U_10U_7_and_9_nl) , m_row0_asn_188 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_12_m1c = ~(IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl = (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_6_else_carry_3_sva);
  assign o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl = nl_o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl[9:0];
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_10_nl = MUX_v_10_2_2((o_col2_3_FpMantRNE_23U_11U_6_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0);
  assign m_row0_and_57_nl = (~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_5) & m_row0_m_row0_nor_12_m1c;
  assign m_row0_and_58_nl = IsNaN_6U_10U_13_land_3_lpi_1_dfm_5 & m_row0_m_row0_nor_12_m1c;
  assign FpAdd_6U_10U_6_o_mant_3_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_10_nl),
      FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_6_o_mant_3_lpi_2,
      {(m_row0_and_57_nl) , (m_row0_and_58_nl) , m_row0_asn_190 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_11_m1c = ~(IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl = (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_6_else_carry_2_sva);
  assign o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl = nl_o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl[9:0];
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_9_nl = MUX_v_10_2_2((o_col2_2_FpMantRNE_23U_11U_6_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0);
  assign m_row0_and_59_nl = (~ IsNaN_6U_10U_13_land_2_lpi_1_dfm_3) & m_row0_m_row0_nor_11_m1c;
  assign m_row0_and_60_nl = IsNaN_6U_10U_13_land_2_lpi_1_dfm_3 & m_row0_m_row0_nor_11_m1c;
  assign FpAdd_6U_10U_6_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_9_nl),
      FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_6_o_mant_2_lpi_2,
      {(m_row0_and_59_nl) , (m_row0_and_60_nl) , m_row0_asn_192 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_10_m1c = ~(IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl = (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_6_else_carry_1_sva);
  assign o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl = nl_o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl[9:0];
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_8_nl = MUX_v_10_2_2((o_col2_1_FpMantRNE_23U_11U_6_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0);
  assign m_row0_and_61_nl = (~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_5) & m_row0_m_row0_nor_10_m1c;
  assign m_row0_and_62_nl = IsNaN_6U_10U_13_land_1_lpi_1_dfm_5 & m_row0_m_row0_nor_10_m1c;
  assign FpAdd_6U_10U_6_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_8_nl),
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_6_o_mant_1_lpi_2,
      {(m_row0_and_61_nl) , (m_row0_and_62_nl) , m_row0_asn_194 , m_row0_unequal_tmp_4});
  assign nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl = FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_2
      + 6'b1;
  assign o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl = nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_31_nl = (~(FpAdd_6U_10U_6_and_2_tmp | FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_19_nl = FpAdd_6U_10U_6_and_2_tmp & (~ FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_32_nl = FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_9_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_21_nl = IsNaN_6U_10U_13_land_3_lpi_1_dfm_5 & (~ IsNaN_6U_10U_11_land_3_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_2,
      (o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_6_o_expo_3_lpi_2,
      {(FpAdd_6U_10U_6_and_31_nl) , (FpAdd_6U_10U_6_and_19_nl) , (FpAdd_6U_10U_6_and_32_nl)
      , (FpAdd_6U_10U_6_and_21_nl) , m_row0_asn_190 , m_row0_unequal_tmp_4});
  assign nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl = FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_2
      + 6'b1;
  assign o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl = nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_29_nl = (~(FpAdd_6U_10U_6_and_1_tmp | FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_13_nl = FpAdd_6U_10U_6_and_1_tmp & (~ FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_30_nl = FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_7_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_15_nl = IsNaN_6U_10U_13_land_2_lpi_1_dfm_3 & (~ IsNaN_6U_10U_11_land_2_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_2,
      (o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_6_o_expo_2_lpi_2,
      {(FpAdd_6U_10U_6_and_29_nl) , (FpAdd_6U_10U_6_and_13_nl) , (FpAdd_6U_10U_6_and_30_nl)
      , (FpAdd_6U_10U_6_and_15_nl) , m_row0_asn_192 , m_row0_unequal_tmp_4});
  assign nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl = FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_2
      + 6'b1;
  assign o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl = nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_nl = (~(FpAdd_6U_10U_6_and_tmp | FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_6_nl = FpAdd_6U_10U_6_and_tmp & (~ FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_28_nl = FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_5_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_9_nl = IsNaN_6U_10U_13_land_1_lpi_1_dfm_5 & (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_2,
      (o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_6_o_expo_1_lpi_2,
      {(FpAdd_6U_10U_6_and_nl) , (FpAdd_6U_10U_6_and_6_nl) , (FpAdd_6U_10U_6_and_28_nl)
      , (FpAdd_6U_10U_6_and_9_nl) , m_row0_asn_194 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_9_m1c = ~(IsNaN_6U_10U_10_land_3_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl = (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_5_else_carry_3_sva);
  assign o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl = nl_o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl[9:0];
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_10_nl = MUX_v_10_2_2((o_col1_3_FpMantRNE_23U_11U_5_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0);
  assign m_row0_and_65_nl = (~ IsNaN_6U_10U_11_land_3_lpi_1_dfm_5) & m_row0_m_row0_nor_9_m1c;
  assign m_row0_and_66_nl = IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 & m_row0_m_row0_nor_9_m1c;
  assign FpAdd_6U_10U_5_o_mant_3_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_10_nl),
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_5_o_mant_3_lpi_2,
      {(m_row0_and_65_nl) , (m_row0_and_66_nl) , m_row0_asn_196 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_8_m1c = ~(IsNaN_6U_10U_10_land_2_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl = (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_5_else_carry_2_sva);
  assign o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl = nl_o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl[9:0];
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_9_nl = MUX_v_10_2_2((o_col1_2_FpMantRNE_23U_11U_5_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0);
  assign m_row0_and_67_nl = (~ IsNaN_6U_10U_11_land_2_lpi_1_dfm_5) & m_row0_m_row0_nor_8_m1c;
  assign m_row0_and_68_nl = IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 & m_row0_m_row0_nor_8_m1c;
  assign FpAdd_6U_10U_5_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_9_nl),
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_5_o_mant_2_lpi_2,
      {(m_row0_and_67_nl) , (m_row0_and_68_nl) , m_row0_asn_198 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_7_m1c = ~(IsNaN_6U_10U_10_land_1_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl = (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_5_else_carry_1_sva);
  assign o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl = nl_o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl[9:0];
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_8_nl = MUX_v_10_2_2((o_col1_1_FpMantRNE_23U_11U_5_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0);
  assign m_row0_and_69_nl = (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_5) & m_row0_m_row0_nor_7_m1c;
  assign m_row0_and_70_nl = IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 & m_row0_m_row0_nor_7_m1c;
  assign FpAdd_6U_10U_5_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_8_nl),
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_5_o_mant_1_lpi_2,
      {(m_row0_and_69_nl) , (m_row0_and_70_nl) , m_row0_asn_200 , m_row0_unequal_tmp_4});
  assign nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl = FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_2
      + 6'b1;
  assign o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl = nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_31_nl = (~(FpAdd_6U_10U_5_and_2_tmp | FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_19_nl = FpAdd_6U_10U_5_and_2_tmp & (~ FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_32_nl = FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_9_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_21_nl = IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 & (~ IsNaN_6U_10U_10_land_3_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_2,
      (o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_5_o_expo_3_lpi_2,
      {(FpAdd_6U_10U_5_and_31_nl) , (FpAdd_6U_10U_5_and_19_nl) , (FpAdd_6U_10U_5_and_32_nl)
      , (FpAdd_6U_10U_5_and_21_nl) , m_row0_asn_196 , m_row0_unequal_tmp_4});
  assign nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl = FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_2
      + 6'b1;
  assign o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl = nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_29_nl = (~(FpAdd_6U_10U_5_and_1_tmp | FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_13_nl = FpAdd_6U_10U_5_and_1_tmp & (~ FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_30_nl = FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_7_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_15_nl = IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 & (~ IsNaN_6U_10U_10_land_2_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_2,
      (o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_5_o_expo_2_lpi_2,
      {(FpAdd_6U_10U_5_and_29_nl) , (FpAdd_6U_10U_5_and_13_nl) , (FpAdd_6U_10U_5_and_30_nl)
      , (FpAdd_6U_10U_5_and_15_nl) , m_row0_asn_198 , m_row0_unequal_tmp_4});
  assign nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl = FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_2
      + 6'b1;
  assign o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl = nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_nl = (~(FpAdd_6U_10U_5_and_tmp | FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_6_nl = FpAdd_6U_10U_5_and_tmp & (~ FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_28_nl = FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_5_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_9_nl = IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 & (~ IsNaN_6U_10U_10_land_1_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_2,
      (o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_5_o_expo_1_lpi_2,
      {(FpAdd_6U_10U_5_and_nl) , (FpAdd_6U_10U_5_and_6_nl) , (FpAdd_6U_10U_5_and_28_nl)
      , (FpAdd_6U_10U_5_and_9_nl) , m_row0_asn_200 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_6_m1c = ~(IsNaN_6U_10U_8_land_3_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl = (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_4_else_carry_3_sva);
  assign o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl = nl_o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl[9:0];
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_10_nl = MUX_v_10_2_2((o_col0_3_FpMantRNE_23U_11U_4_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0);
  assign m_row0_and_73_nl = (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_3) & m_row0_m_row0_nor_6_m1c;
  assign m_row0_and_74_nl = IsNaN_6U_10U_9_land_3_lpi_1_dfm_3 & m_row0_m_row0_nor_6_m1c;
  assign FpAdd_6U_10U_4_o_mant_3_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_10_nl),
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_7, FpAdd_6U_10U_4_o_mant_3_lpi_2,
      {(m_row0_and_73_nl) , (m_row0_and_74_nl) , m_row0_asn_202 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_5_m1c = ~(IsNaN_6U_10U_8_land_2_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl = (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_4_else_carry_2_sva);
  assign o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl = nl_o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl[9:0];
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_9_nl = MUX_v_10_2_2((o_col0_2_FpMantRNE_23U_11U_4_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0);
  assign m_row0_and_75_nl = (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_3) & m_row0_m_row0_nor_5_m1c;
  assign m_row0_and_76_nl = IsNaN_6U_10U_9_land_2_lpi_1_dfm_3 & m_row0_m_row0_nor_5_m1c;
  assign FpAdd_6U_10U_4_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_9_nl),
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_7, FpAdd_6U_10U_4_o_mant_2_lpi_2,
      {(m_row0_and_75_nl) , (m_row0_and_76_nl) , m_row0_asn_204 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_4_m1c = ~(IsNaN_6U_10U_8_land_1_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl = (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_4_else_carry_1_sva);
  assign o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl = nl_o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl[9:0];
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_8_nl = MUX_v_10_2_2((o_col0_1_FpMantRNE_23U_11U_4_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0);
  assign m_row0_and_77_nl = (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_5) & m_row0_m_row0_nor_4_m1c;
  assign m_row0_and_78_nl = IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 & m_row0_m_row0_nor_4_m1c;
  assign FpAdd_6U_10U_4_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_8_nl),
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_o_mant_1_lpi_1_dfm_7, FpAdd_6U_10U_4_o_mant_1_lpi_2,
      {(m_row0_and_77_nl) , (m_row0_and_78_nl) , m_row0_asn_206 , m_row0_unequal_tmp_4});
  assign nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl = FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_2
      + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl = nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_31_nl = (~(FpAdd_6U_10U_4_and_2_tmp | FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_19_nl = FpAdd_6U_10U_4_and_2_tmp & (~ FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_9_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_32_nl = FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_9_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_21_nl = IsNaN_6U_10U_9_land_3_lpi_1_dfm_3 & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_2,
      (o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_4_o_expo_3_lpi_2,
      {(FpAdd_6U_10U_4_and_31_nl) , (FpAdd_6U_10U_4_and_19_nl) , (FpAdd_6U_10U_4_and_32_nl)
      , (FpAdd_6U_10U_4_and_21_nl) , m_row0_asn_202 , m_row0_unequal_tmp_4});
  assign nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl = FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_2
      + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl = nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_29_nl = (~(FpAdd_6U_10U_4_and_1_tmp | FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_13_nl = FpAdd_6U_10U_4_and_1_tmp & (~ FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_7_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_30_nl = FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_7_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_15_nl = IsNaN_6U_10U_9_land_2_lpi_1_dfm_3 & (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_2,
      (o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_4_o_expo_2_lpi_2,
      {(FpAdd_6U_10U_4_and_29_nl) , (FpAdd_6U_10U_4_and_13_nl) , (FpAdd_6U_10U_4_and_30_nl)
      , (FpAdd_6U_10U_4_and_15_nl) , m_row0_asn_204 , m_row0_unequal_tmp_4});
  assign nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl = FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_2
      + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl = nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_nl = (~(FpAdd_6U_10U_4_and_tmp | FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_6_nl = FpAdd_6U_10U_4_and_tmp & (~ FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_5_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_28_nl = FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_5_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_9_nl = IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 & (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_2,
      (o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_4_o_expo_1_lpi_2,
      {(FpAdd_6U_10U_4_and_nl) , (FpAdd_6U_10U_4_and_6_nl) , (FpAdd_6U_10U_4_and_28_nl)
      , (FpAdd_6U_10U_4_and_9_nl) , m_row0_asn_206 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_3_m1c = ~(IsNaN_6U_10U_14_land_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl = (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_7_else_carry_sva);
  assign o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl = nl_o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl[9:0];
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_11_nl = MUX_v_10_2_2((o_col3_4_FpMantRNE_23U_11U_7_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0);
  assign m_row0_and_47_nl = (~ IsNaN_6U_10U_15_land_lpi_1_dfm_5) & m_row0_m_row0_nor_3_m1c;
  assign m_row0_and_48_nl = IsNaN_6U_10U_15_land_lpi_1_dfm_5 & m_row0_m_row0_nor_3_m1c;
  assign FpAdd_6U_10U_7_o_mant_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_7_FpAdd_6U_10U_7_or_11_nl),
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_7, FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_7_o_mant_lpi_2,
      {(m_row0_and_47_nl) , (m_row0_and_48_nl) , m_row0_asn_208 , m_row0_unequal_tmp_4});
  assign nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl = FpAdd_6U_10U_7_o_expo_lpi_1_dfm_2
      + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl = nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_33_nl = (~(FpAdd_6U_10U_7_and_3_tmp | FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_25_nl = FpAdd_6U_10U_7_and_3_tmp & (~ FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_34_nl = FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_11_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_and_27_nl = IsNaN_6U_10U_15_land_lpi_1_dfm_5 & (~ IsNaN_6U_10U_14_land_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_7_o_expo_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_7_o_expo_lpi_1_dfm_2,
      (o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_7_o_expo_lpi_2,
      {(FpAdd_6U_10U_7_and_33_nl) , (FpAdd_6U_10U_7_and_25_nl) , (FpAdd_6U_10U_7_and_34_nl)
      , (FpAdd_6U_10U_7_and_27_nl) , m_row0_asn_208 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_2_m1c = ~(IsNaN_6U_10U_11_land_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl = (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_6_else_carry_sva);
  assign o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl = nl_o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl[9:0];
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_11_nl = MUX_v_10_2_2((o_col2_4_FpMantRNE_23U_11U_6_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0);
  assign m_row0_and_55_nl = (~ IsNaN_6U_10U_13_land_lpi_1_dfm_5) & m_row0_m_row0_nor_2_m1c;
  assign m_row0_and_56_nl = IsNaN_6U_10U_13_land_lpi_1_dfm_5 & m_row0_m_row0_nor_2_m1c;
  assign FpAdd_6U_10U_6_o_mant_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_6_FpAdd_6U_10U_6_or_11_nl),
      FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_6_o_mant_lpi_2,
      {(m_row0_and_55_nl) , (m_row0_and_56_nl) , m_row0_asn_210 , m_row0_unequal_tmp_4});
  assign nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl = FpAdd_6U_10U_6_o_expo_lpi_1_dfm_2
      + 6'b1;
  assign o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl = nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_33_nl = (~(FpAdd_6U_10U_6_and_3_tmp | FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_25_nl = FpAdd_6U_10U_6_and_3_tmp & (~ FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_34_nl = FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_11_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_and_27_nl = IsNaN_6U_10U_13_land_lpi_1_dfm_5 & (~ IsNaN_6U_10U_11_land_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_6_o_expo_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_6_o_expo_lpi_1_dfm_2,
      (o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_6_o_expo_lpi_2,
      {(FpAdd_6U_10U_6_and_33_nl) , (FpAdd_6U_10U_6_and_25_nl) , (FpAdd_6U_10U_6_and_34_nl)
      , (FpAdd_6U_10U_6_and_27_nl) , m_row0_asn_210 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_1_m1c = ~(IsNaN_6U_10U_10_land_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl = (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_5_else_carry_sva);
  assign o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl = nl_o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl[9:0];
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_11_nl = MUX_v_10_2_2((o_col1_4_FpMantRNE_23U_11U_5_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0);
  assign m_row0_and_63_nl = (~ IsNaN_6U_10U_11_land_lpi_1_dfm_5) & m_row0_m_row0_nor_1_m1c;
  assign m_row0_and_64_nl = IsNaN_6U_10U_11_land_lpi_1_dfm_5 & m_row0_m_row0_nor_1_m1c;
  assign FpAdd_6U_10U_5_o_mant_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_5_FpAdd_6U_10U_5_or_11_nl),
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7, FpAdd_6U_10U_5_o_mant_lpi_2,
      {(m_row0_and_63_nl) , (m_row0_and_64_nl) , m_row0_asn_212 , m_row0_unequal_tmp_4});
  assign nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl = FpAdd_6U_10U_5_o_expo_lpi_1_dfm_2
      + 6'b1;
  assign o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl = nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_33_nl = (~(FpAdd_6U_10U_5_and_3_tmp | FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_25_nl = FpAdd_6U_10U_5_and_3_tmp & (~ FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_34_nl = FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_11_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_and_27_nl = IsNaN_6U_10U_11_land_lpi_1_dfm_5 & (~ IsNaN_6U_10U_10_land_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_5_o_expo_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_5_o_expo_lpi_1_dfm_2,
      (o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_5_o_expo_lpi_2,
      {(FpAdd_6U_10U_5_and_33_nl) , (FpAdd_6U_10U_5_and_25_nl) , (FpAdd_6U_10U_5_and_34_nl)
      , (FpAdd_6U_10U_5_and_27_nl) , m_row0_asn_212 , m_row0_unequal_tmp_4});
  assign m_row0_m_row0_nor_m1c = ~(IsNaN_6U_10U_8_land_lpi_1_dfm_5 | m_row0_unequal_tmp_4);
  assign nl_o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl = (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_4_else_carry_sva);
  assign o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl = nl_o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl[9:0];
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_11_nl = MUX_v_10_2_2((o_col0_4_FpMantRNE_23U_11U_4_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0);
  assign m_row0_and_71_nl = (~ IsNaN_6U_10U_9_land_lpi_1_dfm_3) & m_row0_m_row0_nor_m1c;
  assign m_row0_and_72_nl = IsNaN_6U_10U_9_land_lpi_1_dfm_3 & m_row0_m_row0_nor_m1c;
  assign FpAdd_6U_10U_4_o_mant_lpi_1_dfm_3_mx0w0 = MUX1HOT_v_10_4_2((FpAdd_6U_10U_4_FpAdd_6U_10U_4_or_11_nl),
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7, FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_7, FpAdd_6U_10U_4_o_mant_lpi_2,
      {(m_row0_and_71_nl) , (m_row0_and_72_nl) , m_row0_asn_214 , m_row0_unequal_tmp_4});
  assign nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl = FpAdd_6U_10U_4_o_expo_lpi_1_dfm_2
      + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl = nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_33_nl = (~(FpAdd_6U_10U_4_and_3_tmp | FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_25_nl = FpAdd_6U_10U_4_and_3_tmp & (~ FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_11_m1c & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_34_nl = FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_11_m1c
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_and_27_nl = IsNaN_6U_10U_9_land_lpi_1_dfm_3 & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_5)
      & (~ m_row0_unequal_tmp_4);
  assign FpAdd_6U_10U_4_o_expo_lpi_1_dfm_8_mx0w0 = MUX1HOT_v_6_6_2(FpAdd_6U_10U_4_o_expo_lpi_1_dfm_2,
      (o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_nl), 6'b111110, ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2}),
      ({reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_1
      , reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_2}), FpAdd_6U_10U_4_o_expo_lpi_2,
      {(FpAdd_6U_10U_4_and_33_nl) , (FpAdd_6U_10U_4_and_25_nl) , (FpAdd_6U_10U_4_and_34_nl)
      , (FpAdd_6U_10U_4_and_27_nl) , m_row0_asn_214 , m_row0_unequal_tmp_4});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse = IsNaN_6U_10U_7_land_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse;
  assign FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx1 = MUX_v_10_2_2(FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_11_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse = IsNaN_6U_10U_5_land_lpi_1_dfm_3
      | IsNaN_6U_10U_4_land_lpi_1_dfm_st_2;
  assign FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx1 = MUX_v_10_2_2(FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_11_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse = IsNaN_6U_10U_3_land_lpi_1_dfm_3
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_2;
  assign FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx1 = MUX_v_10_2_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_11_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse = IsNaN_6U_10U_1_land_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse;
  assign FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx1 = MUX_v_10_2_2(FpAdd_6U_10U_FpAdd_6U_10U_or_11_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[9:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w4, or_dcpl_69);
  assign m_row2_if_d1_mux_1_cse = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[137:128]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
      or_dcpl_64);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_15_nl
      = (~ (chn_data_in_rsci_d_mxwt[14])) & IsZero_5U_10U_aelse_not_19;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_15_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3 = ({(chn_data_in_rsci_d_mxwt[14])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl)}) | ({{1{IsInf_5U_10U_land_1_lpi_1_dfm}},
      IsInf_5U_10U_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_land_1_lpi_1_dfm}}, IsNaN_5U_10U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[142])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_19}) | ({{1{IsInf_5U_10U_1_land_1_lpi_1_dfm}},
      IsInf_5U_10U_1_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_1_land_1_lpi_1_dfm}},
      IsNaN_5U_10U_1_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[25:16]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_2_mx0w4, or_dcpl_80);
  assign m_row2_if_d1_mux_4_cse = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[153:144]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
      or_dcpl_75);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_14_nl
      = (~ (chn_data_in_rsci_d_mxwt[30])) & IsZero_5U_10U_aelse_not_17;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_14_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3 = ({(chn_data_in_rsci_d_mxwt[30])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl)}) | ({{1{IsInf_5U_10U_land_2_lpi_1_dfm}},
      IsInf_5U_10U_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_land_2_lpi_1_dfm}}, IsNaN_5U_10U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[158])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_21}) | ({{1{IsInf_5U_10U_1_land_2_lpi_1_dfm}},
      IsInf_5U_10U_1_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_1_land_2_lpi_1_dfm}},
      IsNaN_5U_10U_1_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[41:32]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w4, or_dcpl_91);
  assign m_row2_if_d1_mux_7_cse = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[169:160]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
      or_dcpl_86);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_13_nl
      = (~ (chn_data_in_rsci_d_mxwt[46])) & IsZero_5U_10U_aelse_not_15;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_13_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3 = ({(chn_data_in_rsci_d_mxwt[46])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl)}) | ({{1{IsInf_5U_10U_land_3_lpi_1_dfm}},
      IsInf_5U_10U_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_land_3_lpi_1_dfm}}, IsNaN_5U_10U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[174])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_23}) | ({{1{IsInf_5U_10U_1_land_3_lpi_1_dfm}},
      IsInf_5U_10U_1_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_1_land_3_lpi_1_dfm}},
      IsNaN_5U_10U_1_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[73:64]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
      or_dcpl_126);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[78])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_25}) | ({{1{IsInf_5U_10U_2_land_1_lpi_1_dfm}},
      IsInf_5U_10U_2_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_2_land_1_lpi_1_dfm}},
      IsNaN_5U_10U_2_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[89:80]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
      or_dcpl_116);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[94])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_19}) | ({{1{IsInf_5U_10U_2_land_2_lpi_1_dfm}},
      IsInf_5U_10U_2_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_2_land_2_lpi_1_dfm}},
      IsNaN_5U_10U_2_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[105:96]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
      or_dcpl_106);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[110])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_21}) | ({{1{IsInf_5U_10U_2_land_3_lpi_1_dfm}},
      IsInf_5U_10U_2_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_2_land_3_lpi_1_dfm}},
      IsNaN_5U_10U_2_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_1_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[201:192]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_mx0w4,
      or_dcpl_131);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_15_nl
      = (~ (chn_data_in_rsci_d_mxwt[206])) & IsZero_5U_10U_7_aelse_not_19;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_2_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_15_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_7_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[206])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_2_nl)}) | ({{1{IsInf_5U_10U_7_land_1_lpi_1_dfm}},
      IsInf_5U_10U_7_land_1_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_7_land_1_lpi_1_dfm}},
      IsNaN_5U_10U_7_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_2_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[217:208]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_2_mx0w4,
      or_dcpl_121);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_14_nl
      = (~ (chn_data_in_rsci_d_mxwt[222])) & IsZero_5U_10U_7_aelse_not_17;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_7_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_14_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_7_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[222])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_7_nl)}) | ({{1{IsInf_5U_10U_7_land_2_lpi_1_dfm}},
      IsInf_5U_10U_7_land_2_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_7_land_2_lpi_1_dfm}},
      IsNaN_5U_10U_7_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_3_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[233:224]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_4_mx0w4,
      or_dcpl_111);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_13_nl
      = (~ (chn_data_in_rsci_d_mxwt[238])) & IsZero_5U_10U_7_aelse_not_15;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_12_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_13_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_7_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[238])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_12_nl)}) | ({{1{IsInf_5U_10U_7_land_3_lpi_1_dfm}},
      IsInf_5U_10U_7_land_3_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_7_land_3_lpi_1_dfm}},
      IsNaN_5U_10U_7_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_5, or_dcpl_1);
  assign IsZero_5U_10U_1_aelse_not_12_nl = ~ IsZero_5U_10U_1_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_9_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[185:176]), (IsZero_5U_10U_1_aelse_not_12_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_35_nl = MUX_v_10_2_2(m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_9_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux_35_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[57:48]), IsZero_5U_10U_aelse_not_13);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_26_nl = MUX_v_10_2_2(m_row0_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_6_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_26_nl), 10'b1111111111,
      IsInf_5U_10U_land_lpi_1_dfm);
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp = m_row0_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp = m_row0_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp = m_row2_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]) & FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2==4'b1111);
  assign IsZero_5U_10U_2_aelse_not_12_nl = ~ IsZero_5U_10U_2_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_9_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[121:112]), (IsZero_5U_10U_2_aelse_not_12_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_33_nl = MUX_v_10_2_2(m_row1_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_9_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_33_nl), 10'b1111111111,
      IsInf_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_9_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_data_in_rsci_d_mxwt[249:240]), IsZero_5U_10U_7_aelse_not_13);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_27_nl = MUX_v_10_2_2(m_row3_4_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_9_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_6_mx0w4
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux_27_nl), 10'b1111111111,
      IsInf_5U_10U_7_land_lpi_1_dfm);
  assign IsZero_5U_10U_2_aelse_not_20_nl = ~ IsZero_5U_10U_2_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[125:122]), (IsZero_5U_10U_2_aelse_not_20_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_cse
      , IsDenorm_5U_10U_2_land_lpi_1_dfm , IsInf_5U_10U_2_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl),
      4'b1111, IsNaN_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[253:250]), IsZero_5U_10U_7_aelse_not_13);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_3_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_3_cse
      , IsDenorm_5U_10U_7_land_lpi_1_dfm , IsInf_5U_10U_7_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_mux1h_3_nl),
      4'b1111, IsNaN_5U_10U_7_land_lpi_1_dfm);
  assign IsZero_5U_10U_1_aelse_not_20_nl = ~ IsZero_5U_10U_1_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[189:186]), (IsZero_5U_10U_1_aelse_not_20_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_10_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse
      , IsDenorm_5U_10U_1_land_lpi_1_dfm , IsInf_5U_10U_1_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_mux1h_10_nl),
      4'b1111, IsNaN_5U_10U_1_land_lpi_1_dfm);
  assign IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp = m_row2_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3==2'b11) & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2==4'b1111);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_data_in_rsci_d_mxwt[61:58]), IsZero_5U_10U_aelse_not_13);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse
      , IsDenorm_5U_10U_land_lpi_1_dfm , IsInf_5U_10U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl),
      4'b1111, IsNaN_5U_10U_land_lpi_1_dfm);
  assign o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0 = (FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)
      | FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_5 | FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0 = (FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)
      | FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_5 | FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0 = (FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5 | FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0 = (FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)
      | FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5 | FpAdd_6U_10U_o_expo_lpi_1_dfm_7_4 | (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col1_4_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0 = (FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_5 | FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col1_3_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0 = (FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_5 | FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col1_2_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0 = (FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5 | FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col1_1_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0 = (FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5 | FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0 = (FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_5 | FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0 = (FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_5 | FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0 = (FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_5 | FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0 = (FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_5 | FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0 = (FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5 | FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0 = (FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5 | FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0 = (FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5 | FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0!=4'b0000);
  assign o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0 = (FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)
      | FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5 | FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_4
      | (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0!=4'b0000);
  assign data_truncate_equal_tmp_mx0w0 = ~((cfg_precision!=2'b00));
  assign data_truncate_nor_tmp_mx0w0 = ~(((cfg_precision==2'b01)) | data_truncate_equal_tmp_mx0w0);
  assign data_truncate_nor_dfs_mx0w0 = ~(data_truncate_equal_tmp_mx0w0 | data_truncate_nor_tmp_mx0w0);
  assign IsNaN_6U_10U_9_land_2_lpi_1_dfm_mx0w0 = ~(IsNaN_6U_10U_9_nor_1_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm_2);
  assign IsNaN_6U_10U_9_land_3_lpi_1_dfm_mx0w0 = ~(IsNaN_6U_10U_9_nor_2_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm_2);
  assign IsNaN_6U_10U_9_land_lpi_1_dfm_mx0w0 = ~(IsNaN_6U_10U_9_nor_3_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm_2);
  assign IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_2_tmp = ~((~((FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)))
      | (~(FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_5 & FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp = ~((~((FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_5 & FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_1_tmp = ~((~((FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)))
      | (~(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5 & FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp = ~(IsNaN_6U_10U_10_nor_1_tmp
      | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp);
  assign IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_tmp = ~((~((FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)))
      | (~(FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5 & FpAdd_6U_10U_o_expo_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp = ~((~((FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5 & FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp = ~(IsNaN_6U_10U_9_nor_2_tmp |
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp);
  assign IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp = ~(IsNaN_6U_10U_9_nor_1_tmp |
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp);
  assign IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp = ~((~((FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5 & FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp = ~((~((FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_5 & FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp = ~((~((FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5 & FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp = ~((~((FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5 & FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_3_tmp = ~((~((FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx1!=10'b0000000000)))
      | (~(FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_5 & FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp = ~((~((FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_5 & FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_3_0==4'b1111))));
  assign IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp = ~(IsNaN_6U_10U_9_nor_3_tmp |
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp);
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp = ~((~((FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | (~(FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_5 & FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_4
      & (FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_3_0==4'b1111))));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[57:48]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_6_mx0w4, or_dcpl_341);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[185:176]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
      or_dcpl_336);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_12_nl
      = (~ (chn_data_in_rsci_d_mxwt[62])) & IsZero_5U_10U_aelse_not_13;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_12_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3 = ({(chn_data_in_rsci_d_mxwt[62])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl)}) | ({{1{IsInf_5U_10U_land_lpi_1_dfm}},
      IsInf_5U_10U_land_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_land_lpi_1_dfm}}, IsNaN_5U_10U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[190])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_25}) | ({{1{IsInf_5U_10U_1_land_lpi_1_dfm}},
      IsInf_5U_10U_1_land_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_1_land_lpi_1_dfm}}, IsNaN_5U_10U_1_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[121:112]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
      or_dcpl_350);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[126])
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_23}) | ({{1{IsInf_5U_10U_2_land_lpi_1_dfm}},
      IsInf_5U_10U_2_land_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_2_land_lpi_1_dfm}}, IsNaN_5U_10U_2_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5, or_dcpl_1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_mant_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_data_in_rsci_d_mxwt[249:240]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_6_mx0w4,
      or_dcpl_355);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_12_nl
      = (~ (chn_data_in_rsci_d_mxwt[254])) & IsZero_5U_10U_7_aelse_not_13;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_17_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_and_12_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_7_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4 = ({(chn_data_in_rsci_d_mxwt[254])
      , (FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_mux_17_nl)}) | ({{1{IsInf_5U_10U_7_land_lpi_1_dfm}},
      IsInf_5U_10U_7_land_lpi_1_dfm}) | ({{1{IsNaN_5U_10U_7_land_lpi_1_dfm}}, IsNaN_5U_10U_7_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_3_mx0 = MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4,
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_5, or_dcpl_1);
  assign FpAdd_6U_10U_o_sign_or_4_nl = and_dcpl_1131 | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp)
      & and_dcpl_1133);
  assign FpAdd_6U_10U_o_sign_and_3_nl = FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp
      & and_dcpl_1133;
  assign FpAdd_6U_10U_o_sign_mux1h_8_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[15]),
      (~ (chn_data_in_rsci_d_mxwt[143])), (chn_data_in_rsci_d_mxwt[15]), {IsNaN_6U_10U_IsNaN_6U_10U_and_tmp
      , (FpAdd_6U_10U_o_sign_or_4_nl) , (FpAdd_6U_10U_o_sign_and_3_nl)});
  assign o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0
      = (FpAdd_6U_10U_o_sign_mux1h_8_nl) ^ FpAdd_6U_10U_o_sign_3_lpi_1_dfm_1_mx0;
  assign FpAdd_6U_10U_1_o_sign_or_2_nl = and_dcpl_1136 | ((~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp)
      & and_dcpl_1138);
  assign FpAdd_6U_10U_1_o_sign_and_3_nl = FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp
      & and_dcpl_1138;
  assign FpAdd_6U_10U_1_o_sign_mux1h_20_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[79]),
      (chn_data_in_rsci_d_mxwt[143]), (chn_data_in_rsci_d_mxwt[79]), {IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp
      , (FpAdd_6U_10U_1_o_sign_or_2_nl) , (FpAdd_6U_10U_1_o_sign_and_3_nl)});
  assign o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0
      = (FpAdd_6U_10U_1_o_sign_mux1h_20_nl) ^ FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_1_mx0;
  assign m_row1_if_d2_or_4_nl = and_dcpl_1141 | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp)
      & and_dcpl_1143);
  assign m_row1_if_d2_and_3_nl = FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp
      & and_dcpl_1143;
  assign m_row1_if_d2_mux1h_4_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[143]),
      (~ (chn_data_in_rsci_d_mxwt[79])), (chn_data_in_rsci_d_mxwt[143]), {IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp
      , (m_row1_if_d2_or_4_nl) , (m_row1_if_d2_and_3_nl)});
  assign o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0
      = (m_row1_if_d2_mux1h_4_nl) ^ FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_1_mx0;
  assign FpAdd_6U_10U_1_o_sign_or_10_nl = and_dcpl_1146 | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp)
      & and_dcpl_1148);
  assign FpAdd_6U_10U_1_o_sign_and_7_nl = FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp
      & and_dcpl_1148;
  assign FpAdd_6U_10U_1_o_sign_mux1h_24_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[79]),
      (~ (chn_data_in_rsci_d_mxwt[207])), (chn_data_in_rsci_d_mxwt[79]), {IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp
      , (FpAdd_6U_10U_1_o_sign_or_10_nl) , (FpAdd_6U_10U_1_o_sign_and_7_nl)});
  assign o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0
      = (FpAdd_6U_10U_1_o_sign_mux1h_24_nl) ^ FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_1_mx0;
  assign o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0
      = ~(FpAdd_6U_10U_o_sign_2_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_o_sign_3_lpi_1_dfm_1_mx0);
  assign o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0
      = ~(FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_1_mx0);
  assign o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0
      = ~(FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_1_mx0);
  assign o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0
      = ~(FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_1_mx0);
  assign o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_o_sign_3_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_o_sign_2_lpi_1_dfm_1_mx0;
  assign o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_1_mx0;
  assign o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_1_mx0;
  assign o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_1_mx0 ^ FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_1_mx0;
  assign FpAdd_6U_10U_o_sign_or_5_nl = and_dcpl_1206 | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp)
      & and_dcpl_1208);
  assign FpAdd_6U_10U_o_sign_and_7_nl = FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp
      & and_dcpl_1208;
  assign FpAdd_6U_10U_o_sign_mux1h_11_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[63]),
      (~ (chn_data_in_rsci_d_mxwt[191])), (chn_data_in_rsci_d_mxwt[63]), {IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp
      , (FpAdd_6U_10U_o_sign_or_5_nl) , (FpAdd_6U_10U_o_sign_and_7_nl)});
  assign o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_o_sign_2_lpi_1_dfm_1_mx0 ^ (FpAdd_6U_10U_o_sign_mux1h_11_nl);
  assign FpAdd_6U_10U_1_o_sign_or_7_nl = and_dcpl_1201 | ((~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp)
      & and_dcpl_1203);
  assign FpAdd_6U_10U_1_o_sign_and_11_nl = FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp
      & and_dcpl_1203;
  assign FpAdd_6U_10U_1_o_sign_mux1h_23_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[127]),
      (chn_data_in_rsci_d_mxwt[191]), (chn_data_in_rsci_d_mxwt[127]), {IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp
      , (FpAdd_6U_10U_1_o_sign_or_7_nl) , (FpAdd_6U_10U_1_o_sign_and_11_nl)});
  assign o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_1_mx0 ^ (FpAdd_6U_10U_1_o_sign_mux1h_23_nl);
  assign m_row1_if_d2_or_5_nl = and_dcpl_1196 | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp)
      & and_dcpl_1198);
  assign m_row1_if_d2_and_7_nl = FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp
      & and_dcpl_1198;
  assign m_row1_if_d2_mux1h_7_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[191]),
      (~ (chn_data_in_rsci_d_mxwt[127])), (chn_data_in_rsci_d_mxwt[191]), {IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp
      , (m_row1_if_d2_or_5_nl) , (m_row1_if_d2_and_7_nl)});
  assign o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_1_mx0 ^ (m_row1_if_d2_mux1h_7_nl);
  assign FpAdd_6U_10U_1_o_sign_or_11_nl = and_dcpl_1191 | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp)
      & and_dcpl_1193);
  assign FpAdd_6U_10U_1_o_sign_and_15_nl = FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp
      & and_dcpl_1193;
  assign FpAdd_6U_10U_1_o_sign_mux1h_27_nl = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[127]),
      (~ (chn_data_in_rsci_d_mxwt[255])), (chn_data_in_rsci_d_mxwt[127]), {IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp
      , (FpAdd_6U_10U_1_o_sign_or_11_nl) , (FpAdd_6U_10U_1_o_sign_and_15_nl)});
  assign o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0
      = FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_1_mx0 ^ (FpAdd_6U_10U_1_o_sign_mux1h_27_nl);
  assign FpAdd_6U_10U_4_mux_33_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5),
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5, FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1);
  assign FpAdd_6U_10U_4_else_6_mux_6_nl = MUX_s_1_2_2((FpAdd_6U_10U_4_mux_33_nl),
      (~ FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5), IsNaN_6U_10U_9_land_3_lpi_1_dfm_mx0w0);
  assign FpAdd_6U_10U_4_mux_45_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_4_else_6_mux_6_nl),
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5, IsNaN_6U_10U_8_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_4_mux_1_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2),
      FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2, FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1);
  assign FpAdd_6U_10U_4_else_6_mux_nl = MUX_s_1_2_2((FpAdd_6U_10U_4_mux_1_nl), (~
      FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2), IsNaN_6U_10U_12_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_4_mux_13_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_4_else_6_mux_nl),
      FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2, IsNaN_6U_10U_8_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_33_nl = MUX_s_1_2_2(FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5,
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1);
  assign FpAdd_6U_10U_5_else_6_mux_6_nl = MUX_s_1_2_2((FpAdd_6U_10U_5_mux_33_nl),
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_45_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_5_else_6_mux_6_nl),
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_10_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_1_nl = MUX_s_1_2_2(FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2,
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2, FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1);
  assign FpAdd_6U_10U_5_else_6_mux_nl = MUX_s_1_2_2((FpAdd_6U_10U_5_mux_1_nl), FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2,
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_13_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_5_else_6_mux_nl),
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2, IsNaN_6U_10U_10_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_33_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5),
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5, FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1);
  assign FpAdd_6U_10U_6_else_6_mux_6_nl = MUX_s_1_2_2((FpAdd_6U_10U_6_mux_33_nl),
      (~ FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5), IsNaN_6U_10U_13_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_45_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_6_else_6_mux_6_nl),
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_1_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2),
      FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2, FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1);
  assign FpAdd_6U_10U_6_else_6_mux_nl = MUX_s_1_2_2((FpAdd_6U_10U_6_mux_1_nl), (~
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2), IsNaN_6U_10U_13_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_13_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_6_else_6_mux_nl),
      FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2, IsNaN_6U_10U_12_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_4_mux_17_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5),
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5, FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1);
  assign FpAdd_6U_10U_4_else_6_mux_3_nl = MUX_s_1_2_2((FpAdd_6U_10U_4_mux_17_nl),
      (~ FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5), IsNaN_6U_10U_9_land_2_lpi_1_dfm_mx0w0);
  assign FpAdd_6U_10U_4_mux_29_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_4_else_6_mux_3_nl),
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5, IsNaN_6U_10U_8_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_17_nl = MUX_s_1_2_2(FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5,
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1);
  assign FpAdd_6U_10U_5_else_6_mux_3_nl = MUX_s_1_2_2((FpAdd_6U_10U_5_mux_17_nl),
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_29_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_5_else_6_mux_3_nl),
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_10_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_17_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5),
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5, FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1);
  assign FpAdd_6U_10U_6_else_6_mux_3_nl = MUX_s_1_2_2((FpAdd_6U_10U_6_mux_17_nl),
      (~ FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5), nor_384_cse);
  assign FpAdd_6U_10U_6_mux_29_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_6_else_6_mux_3_nl),
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_4_mux_49_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5),
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5, FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1);
  assign FpAdd_6U_10U_4_else_6_mux_9_nl = MUX_s_1_2_2((FpAdd_6U_10U_4_mux_49_nl),
      (~ FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5), IsNaN_6U_10U_9_land_lpi_1_dfm_mx0w0);
  assign FpAdd_6U_10U_4_mux_61_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_4_else_6_mux_9_nl),
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5, IsNaN_6U_10U_8_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_49_nl = MUX_s_1_2_2(FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5,
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1);
  assign FpAdd_6U_10U_5_else_6_mux_9_nl = MUX_s_1_2_2((FpAdd_6U_10U_5_mux_49_nl),
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_5_mux_61_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_5_else_6_mux_9_nl),
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_10_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_49_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5),
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5, FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1);
  assign FpAdd_6U_10U_6_else_6_mux_9_nl = MUX_s_1_2_2((FpAdd_6U_10U_6_mux_49_nl),
      (~ FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5), IsNaN_6U_10U_13_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_6_mux_61_mx1w1 = MUX_s_1_2_2((FpAdd_6U_10U_6_else_6_mux_9_nl),
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5, IsNaN_6U_10U_12_land_lpi_1_dfm_4);
  assign IsNaN_6U_10U_9_nor_1_tmp = ~((FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000));
  assign IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp = ~(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5
      & FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4 & (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0==4'b1111));
  assign IsNaN_6U_10U_9_nor_2_tmp = ~((FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000));
  assign IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp = ~(FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_5
      & FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_4 & (FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0==4'b1111));
  assign IsNaN_6U_10U_9_nor_3_tmp = ~((FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000));
  assign IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp = ~(FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_5
      & FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_4 & (FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_3_0==4'b1111));
  assign data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[20]));
  assign data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[20]));
  assign data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[20]));
  assign data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[20]));
  assign data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[20]));
  assign data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[20]));
  assign data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[20]));
  assign data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[20]));
  assign data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[20]));
  assign data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[20]));
  assign data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[20]));
  assign data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[20]));
  assign data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[20]));
  assign data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[20]));
  assign data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[20]));
  assign data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0 = (IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[0])
      | (IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[1]) | (~ (IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[20]));
  assign FpAdd_6U_10U_7_mux_1_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2),
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2, FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1);
  assign FpAdd_6U_10U_7_else_6_mux_nl = MUX_s_1_2_2((FpAdd_6U_10U_7_mux_1_nl), (~
      FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2), IsNaN_6U_10U_15_land_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_7_mux_13_mx1w0 = MUX_s_1_2_2((FpAdd_6U_10U_7_else_6_mux_nl),
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2, IsNaN_6U_10U_14_land_1_lpi_1_dfm_st);
  assign FpAdd_6U_10U_7_mux_17_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5),
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1);
  assign FpAdd_6U_10U_7_else_6_mux_3_nl = MUX_s_1_2_2((FpAdd_6U_10U_7_mux_17_nl),
      (~ FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5), IsNaN_6U_10U_15_land_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_7_mux_29_mx1w0 = MUX_s_1_2_2((FpAdd_6U_10U_7_else_6_mux_3_nl),
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_14_land_2_lpi_1_dfm_st);
  assign FpAdd_6U_10U_7_mux_33_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5),
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1);
  assign FpAdd_6U_10U_7_else_6_mux_6_nl = MUX_s_1_2_2((FpAdd_6U_10U_7_mux_33_nl),
      (~ FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5), IsNaN_6U_10U_15_land_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_7_mux_45_mx1w0 = MUX_s_1_2_2((FpAdd_6U_10U_7_else_6_mux_6_nl),
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_14_land_3_lpi_1_dfm_st);
  assign FpAdd_6U_10U_7_mux_49_nl = MUX_s_1_2_2((~ FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5),
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5, FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1);
  assign FpAdd_6U_10U_7_else_6_mux_9_nl = MUX_s_1_2_2((FpAdd_6U_10U_7_mux_49_nl),
      (~ FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5), IsNaN_6U_10U_15_land_lpi_1_dfm_4);
  assign FpAdd_6U_10U_7_mux_61_mx1w0 = MUX_s_1_2_2((FpAdd_6U_10U_7_else_6_mux_9_nl),
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5, IsNaN_6U_10U_14_land_lpi_1_dfm_st);
  assign FpAdd_6U_10U_1_mux_19_mx0w2 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[159]),
      (chn_data_in_rsci_d_mxwt[95]), FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp);
  assign FpAdd_6U_10U_1_mux_36_mx0w2 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[175]),
      (chn_data_in_rsci_d_mxwt[111]), FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp);
  assign nl_IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[255:240])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[127:112]);
  assign IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0[16:0];
  assign nl_m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[95:80])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[223:208]);
  assign m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0 = nl_m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[127:112])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[191:176]);
  assign IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0[16:0];
  assign nl_m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[159:144])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[95:80]);
  assign m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0 = nl_m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0 = conv_s2s_16_17(~ (chn_data_in_rsci_d_mxwt[127:112]))
      + conv_s2s_16_17(~ (chn_data_in_rsci_d_mxwt[191:176])) + 17'b1;
  assign IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0 = nl_IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0[16:0];
  assign nl_m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[95:80])
      + conv_s2s_16_17(chn_data_in_rsci_d_mxwt[159:144]);
  assign m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = nl_m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[191:176])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[63:48]);
  assign IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0[16:0];
  assign nl_m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[31:16])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[159:144]);
  assign m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = nl_m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[111:96])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[239:224]);
  assign m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0 = nl_m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[175:160])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[111:96]);
  assign m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0 = nl_m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[111:96])
      + conv_s2s_16_17(chn_data_in_rsci_d_mxwt[175:160]);
  assign m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = nl_m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[47:32])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[175:160]);
  assign m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0 = nl_m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0[16:0];
  assign nl_IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[79:64])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[207:192]);
  assign IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0[16:0];
  assign nl_IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[143:128])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[79:64]);
  assign IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0[16:0];
  assign nl_IntAddExt_16U_16U_17U_o_acc_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[79:64])
      + conv_s2s_16_17(chn_data_in_rsci_d_mxwt[143:128]) + 17'b1;
  assign IntAddExt_16U_16U_17U_o_acc_itm_mx0w0 = nl_IntAddExt_16U_16U_17U_o_acc_itm_mx0w0[16:0];
  assign nl_IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0 = conv_s2s_16_17(chn_data_in_rsci_d_mxwt[15:0])
      - conv_s2s_16_17(chn_data_in_rsci_d_mxwt[143:128]);
  assign IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0 = nl_IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0[16:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_32)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_33)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_34)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_35)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_36)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_37)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_38)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_39)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_40)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_19 | IsInf_5U_10U_1_land_1_lpi_1_dfm
      | IsNaN_5U_10U_1_land_1_lpi_1_dfm;
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_41)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_21 | IsInf_5U_10U_1_land_2_lpi_1_dfm
      | IsNaN_5U_10U_1_land_2_lpi_1_dfm;
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_42)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_23 | IsInf_5U_10U_1_land_3_lpi_1_dfm
      | IsNaN_5U_10U_1_land_3_lpi_1_dfm;
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_43)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_25 | IsInf_5U_10U_1_land_lpi_1_dfm
      | IsNaN_5U_10U_1_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_25 | IsInf_5U_10U_2_land_1_lpi_1_dfm
      | IsNaN_5U_10U_2_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_19 | IsInf_5U_10U_2_land_2_lpi_1_dfm
      | IsNaN_5U_10U_2_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_21 | IsInf_5U_10U_2_land_3_lpi_1_dfm
      | IsNaN_5U_10U_2_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      = FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_23 | IsInf_5U_10U_2_land_lpi_1_dfm
      | IsNaN_5U_10U_2_land_lpi_1_dfm;
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_44)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_1_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_45)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_2_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_46)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_3_sva[4:0];
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_811c7f8d09c77d8c18ba8b9e2492b26a3d5a_47)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_7_if_1_if_acc_psp_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_3_cse
      = ~(IsDenorm_5U_10U_7_land_lpi_1_dfm | IsInf_5U_10U_7_land_lpi_1_dfm);
  assign IsDenorm_5U_10U_7_land_lpi_1_dfm = IsDenorm_5U_10U_7_or_3_tmp & IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_sva;
  assign IsInf_5U_10U_7_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[249:240]!=10'b0000000000)
      | (~ IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_sva));
  assign IsNaN_5U_10U_7_land_lpi_1_dfm = IsDenorm_5U_10U_7_or_3_tmp & IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_sva;
  assign IsDenorm_5U_10U_7_or_3_tmp = (chn_data_in_rsci_d_mxwt[249:240]!=10'b0000000000);
  assign IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_sva = (chn_data_in_rsci_d_mxwt[254:250]==5'b11111);
  assign IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_sva = ~((chn_data_in_rsci_d_mxwt[254:250]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_cse
      = ~(IsDenorm_5U_10U_2_land_lpi_1_dfm | IsInf_5U_10U_2_land_lpi_1_dfm);
  assign IsInf_5U_10U_2_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[121:112]!=10'b0000000000)
      | (~ IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_sva));
  assign IsNaN_5U_10U_2_land_lpi_1_dfm = IsDenorm_5U_10U_2_or_3_tmp & IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_sva;
  assign IsDenorm_5U_10U_2_land_lpi_1_dfm = IsDenorm_5U_10U_2_or_3_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_2_cse
      = ~(IsDenorm_5U_10U_7_land_3_lpi_1_dfm | IsInf_5U_10U_7_land_3_lpi_1_dfm);
  assign IsDenorm_5U_10U_7_land_3_lpi_1_dfm = IsDenorm_5U_10U_7_or_2_tmp & IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_3_sva;
  assign IsInf_5U_10U_7_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[233:224]!=10'b0000000000)
      | (~ IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_3_sva));
  assign IsNaN_5U_10U_7_land_3_lpi_1_dfm = IsDenorm_5U_10U_7_or_2_tmp & IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_3_sva;
  assign IsDenorm_5U_10U_7_or_2_tmp = (chn_data_in_rsci_d_mxwt[233:224]!=10'b0000000000);
  assign IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_3_sva = (chn_data_in_rsci_d_mxwt[238:234]==5'b11111);
  assign IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_3_sva = ~((chn_data_in_rsci_d_mxwt[238:234]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_cse
      = ~(IsDenorm_5U_10U_2_land_3_lpi_1_dfm | IsInf_5U_10U_2_land_3_lpi_1_dfm);
  assign IsInf_5U_10U_2_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[105:96]!=10'b0000000000)
      | (~ IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_3_sva));
  assign IsNaN_5U_10U_2_land_3_lpi_1_dfm = IsDenorm_5U_10U_2_or_2_tmp & IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_3_sva;
  assign IsDenorm_5U_10U_2_land_3_lpi_1_dfm = IsDenorm_5U_10U_2_or_2_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_1_cse
      = ~(IsDenorm_5U_10U_7_land_2_lpi_1_dfm | IsInf_5U_10U_7_land_2_lpi_1_dfm);
  assign IsDenorm_5U_10U_7_land_2_lpi_1_dfm = IsDenorm_5U_10U_7_or_1_tmp & IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_2_sva;
  assign IsInf_5U_10U_7_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[217:208]!=10'b0000000000)
      | (~ IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_2_sva));
  assign IsNaN_5U_10U_7_land_2_lpi_1_dfm = IsDenorm_5U_10U_7_or_1_tmp & IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_2_sva;
  assign IsDenorm_5U_10U_7_or_1_tmp = (chn_data_in_rsci_d_mxwt[217:208]!=10'b0000000000);
  assign IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_2_sva = (chn_data_in_rsci_d_mxwt[222:218]==5'b11111);
  assign IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_2_sva = ~((chn_data_in_rsci_d_mxwt[222:218]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_cse
      = ~(IsDenorm_5U_10U_2_land_2_lpi_1_dfm | IsInf_5U_10U_2_land_2_lpi_1_dfm);
  assign IsInf_5U_10U_2_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[89:80]!=10'b0000000000)
      | (~ IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_2_sva));
  assign IsNaN_5U_10U_2_land_2_lpi_1_dfm = IsDenorm_5U_10U_2_or_1_tmp & IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_2_sva;
  assign IsDenorm_5U_10U_2_land_2_lpi_1_dfm = IsDenorm_5U_10U_2_or_1_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_nor_cse
      = ~(IsDenorm_5U_10U_7_land_1_lpi_1_dfm | IsInf_5U_10U_7_land_1_lpi_1_dfm);
  assign IsDenorm_5U_10U_7_land_1_lpi_1_dfm = IsDenorm_5U_10U_7_or_tmp & IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_1_sva;
  assign IsInf_5U_10U_7_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[201:192]!=10'b0000000000)
      | (~ IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_1_sva));
  assign IsNaN_5U_10U_7_land_1_lpi_1_dfm = IsDenorm_5U_10U_7_or_tmp & IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_1_sva;
  assign IsDenorm_5U_10U_7_or_tmp = (chn_data_in_rsci_d_mxwt[201:192]!=10'b0000000000);
  assign IsInf_5U_10U_7_IsInf_5U_10U_7_and_cse_1_sva = (chn_data_in_rsci_d_mxwt[206:202]==5'b11111);
  assign IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_1_sva = ~((chn_data_in_rsci_d_mxwt[206:202]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_cse
      = ~(IsDenorm_5U_10U_2_land_1_lpi_1_dfm | IsInf_5U_10U_2_land_1_lpi_1_dfm);
  assign IsInf_5U_10U_2_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[73:64]!=10'b0000000000)
      | (~ IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_1_sva));
  assign IsNaN_5U_10U_2_land_1_lpi_1_dfm = IsDenorm_5U_10U_2_or_tmp & IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_1_sva;
  assign IsDenorm_5U_10U_2_land_1_lpi_1_dfm = IsDenorm_5U_10U_2_or_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse
      = ~(IsDenorm_5U_10U_1_land_lpi_1_dfm | IsInf_5U_10U_1_land_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[185:176]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva));
  assign IsNaN_5U_10U_1_land_lpi_1_dfm = IsDenorm_5U_10U_1_or_3_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva;
  assign IsDenorm_5U_10U_1_land_lpi_1_dfm = IsDenorm_5U_10U_1_or_3_tmp & IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse
      = ~(IsDenorm_5U_10U_1_land_3_lpi_1_dfm | IsInf_5U_10U_1_land_3_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[169:160]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva));
  assign IsNaN_5U_10U_1_land_3_lpi_1_dfm = IsDenorm_5U_10U_1_or_2_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva;
  assign IsDenorm_5U_10U_1_land_3_lpi_1_dfm = IsDenorm_5U_10U_1_or_2_tmp & IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_3_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse
      = ~(IsDenorm_5U_10U_1_land_2_lpi_1_dfm | IsInf_5U_10U_1_land_2_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[153:144]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva));
  assign IsNaN_5U_10U_1_land_2_lpi_1_dfm = IsDenorm_5U_10U_1_or_1_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva;
  assign IsDenorm_5U_10U_1_land_2_lpi_1_dfm = IsDenorm_5U_10U_1_or_1_tmp & IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_2_sva;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse
      = ~(IsDenorm_5U_10U_1_land_1_lpi_1_dfm | IsInf_5U_10U_1_land_1_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[137:128]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva));
  assign IsNaN_5U_10U_1_land_1_lpi_1_dfm = IsDenorm_5U_10U_1_or_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva;
  assign IsDenorm_5U_10U_1_land_1_lpi_1_dfm = IsDenorm_5U_10U_1_or_tmp & IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_1_sva;
  assign IsZero_5U_10U_2_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[121:112]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva));
  assign IsDenorm_5U_10U_2_or_3_tmp = (chn_data_in_rsci_d_mxwt[121:112]!=10'b0000000000);
  assign IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_sva = (chn_data_in_rsci_d_mxwt[126:122]==5'b11111);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva = ~((chn_data_in_rsci_d_mxwt[126:122]!=5'b00000));
  assign IsZero_5U_10U_2_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[105:96]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva));
  assign IsDenorm_5U_10U_2_or_2_tmp = (chn_data_in_rsci_d_mxwt[105:96]!=10'b0000000000);
  assign IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_3_sva = (chn_data_in_rsci_d_mxwt[110:106]==5'b11111);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva = ~((chn_data_in_rsci_d_mxwt[110:106]!=5'b00000));
  assign IsZero_5U_10U_2_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[89:80]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva));
  assign IsDenorm_5U_10U_2_or_1_tmp = (chn_data_in_rsci_d_mxwt[89:80]!=10'b0000000000);
  assign IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_2_sva = (chn_data_in_rsci_d_mxwt[94:90]==5'b11111);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva = ~((chn_data_in_rsci_d_mxwt[94:90]!=5'b00000));
  assign IsZero_5U_10U_2_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[73:64]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva));
  assign IsDenorm_5U_10U_2_or_tmp = (chn_data_in_rsci_d_mxwt[73:64]!=10'b0000000000);
  assign IsInf_5U_10U_2_IsInf_5U_10U_2_and_cse_1_sva = (chn_data_in_rsci_d_mxwt[78:74]==5'b11111);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva = ~((chn_data_in_rsci_d_mxwt[78:74]!=5'b00000));
  assign IsZero_5U_10U_1_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[185:176]!=10'b0000000000)
      | (~ IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_sva));
  assign IsDenorm_5U_10U_1_or_3_tmp = (chn_data_in_rsci_d_mxwt[185:176]!=10'b0000000000);
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva = (chn_data_in_rsci_d_mxwt[190:186]==5'b11111);
  assign IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_sva = ~((chn_data_in_rsci_d_mxwt[190:186]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse
      = ~(IsDenorm_5U_10U_land_lpi_1_dfm | IsInf_5U_10U_land_lpi_1_dfm);
  assign IsDenorm_5U_10U_land_lpi_1_dfm = IsDenorm_5U_10U_or_3_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva;
  assign IsInf_5U_10U_land_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[57:48]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_sva));
  assign IsNaN_5U_10U_land_lpi_1_dfm = IsDenorm_5U_10U_or_3_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_sva;
  assign IsDenorm_5U_10U_or_3_tmp = (chn_data_in_rsci_d_mxwt[57:48]!=10'b0000000000);
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_sva = (chn_data_in_rsci_d_mxwt[62:58]==5'b11111);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva = ~((chn_data_in_rsci_d_mxwt[62:58]!=5'b00000));
  assign IsZero_5U_10U_1_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[169:160]!=10'b0000000000)
      | (~ IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_3_sva));
  assign IsDenorm_5U_10U_1_or_2_tmp = (chn_data_in_rsci_d_mxwt[169:160]!=10'b0000000000);
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva = (chn_data_in_rsci_d_mxwt[174:170]==5'b11111);
  assign IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_3_sva = ~((chn_data_in_rsci_d_mxwt[174:170]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse
      = ~(IsDenorm_5U_10U_land_3_lpi_1_dfm | IsInf_5U_10U_land_3_lpi_1_dfm);
  assign IsDenorm_5U_10U_land_3_lpi_1_dfm = IsDenorm_5U_10U_or_2_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva;
  assign IsInf_5U_10U_land_3_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[41:32]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva));
  assign IsNaN_5U_10U_land_3_lpi_1_dfm = IsDenorm_5U_10U_or_2_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva;
  assign IsDenorm_5U_10U_or_2_tmp = (chn_data_in_rsci_d_mxwt[41:32]!=10'b0000000000);
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva = (chn_data_in_rsci_d_mxwt[46:42]==5'b11111);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva = ~((chn_data_in_rsci_d_mxwt[46:42]!=5'b00000));
  assign IsZero_5U_10U_1_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[153:144]!=10'b0000000000)
      | (~ IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_2_sva));
  assign IsDenorm_5U_10U_1_or_1_tmp = (chn_data_in_rsci_d_mxwt[153:144]!=10'b0000000000);
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva = (chn_data_in_rsci_d_mxwt[158:154]==5'b11111);
  assign IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_2_sva = ~((chn_data_in_rsci_d_mxwt[158:154]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse
      = ~(IsDenorm_5U_10U_land_2_lpi_1_dfm | IsInf_5U_10U_land_2_lpi_1_dfm);
  assign IsDenorm_5U_10U_land_2_lpi_1_dfm = IsDenorm_5U_10U_or_1_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva;
  assign IsInf_5U_10U_land_2_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[25:16]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva));
  assign IsNaN_5U_10U_land_2_lpi_1_dfm = IsDenorm_5U_10U_or_1_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva;
  assign IsDenorm_5U_10U_or_1_tmp = (chn_data_in_rsci_d_mxwt[25:16]!=10'b0000000000);
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva = (chn_data_in_rsci_d_mxwt[30:26]==5'b11111);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva = ~((chn_data_in_rsci_d_mxwt[30:26]!=5'b00000));
  assign IsZero_5U_10U_1_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[137:128]!=10'b0000000000)
      | (~ IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_1_sva));
  assign IsDenorm_5U_10U_1_or_tmp = (chn_data_in_rsci_d_mxwt[137:128]!=10'b0000000000);
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva = (chn_data_in_rsci_d_mxwt[142:138]==5'b11111);
  assign IsZero_5U_10U_1_IsZero_5U_10U_1_nor_cse_1_sva = ~((chn_data_in_rsci_d_mxwt[142:138]!=5'b00000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse =
      ~(IsDenorm_5U_10U_land_1_lpi_1_dfm | IsInf_5U_10U_land_1_lpi_1_dfm);
  assign IsDenorm_5U_10U_land_1_lpi_1_dfm = IsDenorm_5U_10U_or_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva;
  assign IsInf_5U_10U_land_1_lpi_1_dfm = ~((chn_data_in_rsci_d_mxwt[9:0]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva));
  assign IsNaN_5U_10U_land_1_lpi_1_dfm = IsDenorm_5U_10U_or_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva;
  assign IsDenorm_5U_10U_or_tmp = (chn_data_in_rsci_d_mxwt[9:0]!=10'b0000000000);
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva = (chn_data_in_rsci_d_mxwt[14:10]==5'b11111);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva = ~((chn_data_in_rsci_d_mxwt[14:10]!=5'b00000));
  assign nl_FpAdd_6U_10U_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_1_sva = nl_FpAdd_6U_10U_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2, FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_int_mant_p1_1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_int_mant_p1_1_sva_1 = nl_FpAdd_6U_10U_int_mant_p1_1_sva_1[23:0];
  assign FpAdd_6U_10U_o_expo_mux_11_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_o_expo_1_sva_1[5]), m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_o_expo_mux_11_nl), FpAdd_6U_10U_mux_3_itm);
  assign FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_nl = ~(m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_mux_3_itm));
  assign FpAdd_6U_10U_o_expo_and_7_nl = m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_mux_3_itm;
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3,
      (FpAdd_6U_10U_o_expo_1_sva_1[3:0]), (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_nl) , (FpAdd_6U_10U_o_expo_and_7_nl)
      , (~ FpAdd_6U_10U_mux_3_itm)});
  assign FpAdd_6U_10U_o_expo_mux_13_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_o_expo_1_sva_1[4]), m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_o_expo_mux_13_nl), FpAdd_6U_10U_mux_3_itm);
  assign nl_m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_mux_3_itm);
  assign FpMantRNE_23U_11U_else_carry_1_sva = (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_o_expo_1_sva_1 = ({reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_1_sva_1 = nl_FpAdd_6U_10U_o_expo_1_sva_1[5:0];
  assign FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row0_1_FpNormalize_6U_23U_else_lshift_itm, FpNormalize_6U_23U_oelse_not_9);
  assign FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_int_mant_p1_1_sva_1[22:0]),
      (FpAdd_6U_10U_int_mant_p1_1_sva[22:0]), reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_1_sva_1,
      FpAdd_6U_10U_int_mant_p1_1_sva, reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign nl_m_row0_1_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_32)})
      + 6'b1;
  assign m_row0_1_FpNormalize_6U_23U_else_acc_nl = nl_m_row0_1_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row0_1_FpNormalize_6U_23U_else_acc_nl),
      FpNormalize_6U_23U_oelse_not_9);
  assign nl_FpAdd_6U_10U_o_expo_1_sva_4 = ({FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_1_sva_4 = nl_FpAdd_6U_10U_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl = FpAdd_6U_10U_is_inf_1_lpi_1_dfm
      | (~ m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl), m_row0_1_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_is_inf_1_lpi_1_dfm = ~(m_row0_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1[23])));
  assign nl_m_row0_1_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_1_sva);
  assign m_row0_1_FpMantRNE_23U_11U_else_acc_nl = nl_m_row0_1_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_4_itm = MUX_v_10_2_2((m_row0_1_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_2_sva = nl_FpAdd_6U_10U_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2, FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_int_mant_p1_2_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_int_mant_p1_2_sva_1 = nl_FpAdd_6U_10U_int_mant_p1_2_sva_1[23:0];
  assign FpAdd_6U_10U_o_expo_mux_17_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_o_expo_2_sva_1[5]), m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_o_expo_mux_17_nl), FpAdd_6U_10U_mux_20_itm);
  assign FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_1_nl = ~(m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_mux_20_itm));
  assign FpAdd_6U_10U_o_expo_and_5_nl = m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_mux_20_itm;
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3,
      (FpAdd_6U_10U_o_expo_2_sva_1[3:0]), (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_1_nl) , (FpAdd_6U_10U_o_expo_and_5_nl)
      , (~ FpAdd_6U_10U_mux_20_itm)});
  assign FpAdd_6U_10U_o_expo_mux_19_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_o_expo_2_sva_1[4]), m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_o_expo_mux_19_nl), FpAdd_6U_10U_mux_20_itm);
  assign nl_m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_mux_20_itm);
  assign FpMantRNE_23U_11U_else_carry_2_sva = (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_o_expo_2_sva_1 = ({reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_2_sva_1 = nl_FpAdd_6U_10U_o_expo_2_sva_1[5:0];
  assign FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row0_2_FpNormalize_6U_23U_else_lshift_itm, FpNormalize_6U_23U_oelse_not_11);
  assign FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_int_mant_p1_2_sva_1[22:0]),
      (FpAdd_6U_10U_int_mant_p1_2_sva[22:0]), reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_2_sva_1,
      FpAdd_6U_10U_int_mant_p1_2_sva, reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign nl_m_row0_2_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_33)})
      + 6'b1;
  assign m_row0_2_FpNormalize_6U_23U_else_acc_nl = nl_m_row0_2_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row0_2_FpNormalize_6U_23U_else_acc_nl),
      FpNormalize_6U_23U_oelse_not_11);
  assign nl_FpAdd_6U_10U_o_expo_2_sva_4 = ({FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_2_sva_4 = nl_FpAdd_6U_10U_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl = FpAdd_6U_10U_is_inf_2_lpi_1_dfm
      | (~ m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl), m_row0_2_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_is_inf_2_lpi_1_dfm = ~(m_row0_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1[23])));
  assign nl_m_row0_2_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_2_sva);
  assign m_row0_2_FpMantRNE_23U_11U_else_acc_nl = nl_m_row0_2_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_5_itm = MUX_v_10_2_2((m_row0_2_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_3_sva = nl_FpAdd_6U_10U_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2, FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_int_mant_p1_3_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_int_mant_p1_3_sva_1 = nl_FpAdd_6U_10U_int_mant_p1_3_sva_1[23:0];
  assign FpAdd_6U_10U_o_expo_mux_23_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_o_expo_3_sva_1[5]), m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_o_expo_mux_23_nl), FpAdd_6U_10U_mux_37_itm);
  assign FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_2_nl = ~(m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_mux_37_itm));
  assign FpAdd_6U_10U_o_expo_and_3_nl = m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_mux_37_itm;
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3,
      (FpAdd_6U_10U_o_expo_3_sva_1[3:0]), (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_2_nl) , (FpAdd_6U_10U_o_expo_and_3_nl)
      , (~ FpAdd_6U_10U_mux_37_itm)});
  assign FpAdd_6U_10U_o_expo_mux_25_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_o_expo_3_sva_1[4]), m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_o_expo_mux_25_nl), FpAdd_6U_10U_mux_37_itm);
  assign nl_m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_mux_37_itm);
  assign FpMantRNE_23U_11U_else_carry_3_sva = (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_o_expo_3_sva_1 = ({reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_3_sva_1 = nl_FpAdd_6U_10U_o_expo_3_sva_1[5:0];
  assign FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row0_3_FpNormalize_6U_23U_else_lshift_itm, FpNormalize_6U_23U_oelse_not_13);
  assign FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_int_mant_p1_3_sva_1[22:0]),
      (FpAdd_6U_10U_int_mant_p1_3_sva[22:0]), reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_3_sva_1,
      FpAdd_6U_10U_int_mant_p1_3_sva, reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign nl_m_row0_3_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_34)})
      + 6'b1;
  assign m_row0_3_FpNormalize_6U_23U_else_acc_nl = nl_m_row0_3_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row0_3_FpNormalize_6U_23U_else_acc_nl),
      FpNormalize_6U_23U_oelse_not_13);
  assign nl_FpAdd_6U_10U_o_expo_3_sva_4 = ({FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_3_sva_4 = nl_FpAdd_6U_10U_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl = FpAdd_6U_10U_is_inf_3_lpi_1_dfm
      | (~ m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl), m_row0_3_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_is_inf_3_lpi_1_dfm = ~(m_row0_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1[23])));
  assign nl_m_row0_3_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_3_sva);
  assign m_row0_3_FpMantRNE_23U_11U_else_acc_nl = nl_m_row0_3_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_6_itm = MUX_v_10_2_2((m_row0_3_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_sva = nl_FpAdd_6U_10U_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_sva_2, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_sva_2, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_int_mant_p1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_int_mant_p1_sva_1 = nl_FpAdd_6U_10U_int_mant_p1_sva_1[23:0];
  assign FpAdd_6U_10U_o_expo_mux_29_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_o_expo_sva_1[5]), m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_o_expo_mux_29_nl), FpAdd_6U_10U_mux_69_itm);
  assign FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_3_nl = ~(m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_mux_69_itm));
  assign FpAdd_6U_10U_o_expo_and_1_nl = m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_mux_69_itm;
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3,
      (FpAdd_6U_10U_o_expo_sva_1[3:0]), (FpAdd_6U_10U_o_expo_lpi_1_dfm_1[3:0]), {(FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_3_nl)
      , (FpAdd_6U_10U_o_expo_and_1_nl) , (~ FpAdd_6U_10U_mux_69_itm)});
  assign FpAdd_6U_10U_o_expo_mux_31_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_o_expo_sva_1[4]), m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_o_expo_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_o_expo_mux_31_nl), FpAdd_6U_10U_mux_69_itm);
  assign nl_FpAdd_6U_10U_o_expo_sva_1 = ({reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_sva_1 = nl_FpAdd_6U_10U_o_expo_sva_1[5:0];
  assign nl_m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row0_4_FpNormalize_6U_23U_else_lshift_itm, FpNormalize_6U_23U_oelse_not_15);
  assign FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_int_mant_p1_sva_1[22:0]),
      (FpAdd_6U_10U_int_mant_p1_sva[22:0]), reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_sva_1,
      FpAdd_6U_10U_int_mant_p1_sva, reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign nl_m_row0_4_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_35)})
      + 6'b1;
  assign m_row0_4_FpNormalize_6U_23U_else_acc_nl = nl_m_row0_4_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row0_4_FpNormalize_6U_23U_else_acc_nl),
      FpNormalize_6U_23U_oelse_not_15);
  assign nl_m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_o_expo_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_1_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_1_sva = nl_FpAdd_6U_10U_1_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_1_a_int_mant_p1_1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_1_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1[23:0];
  assign FpAdd_6U_10U_1_o_expo_mux_11_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_1_o_expo_1_sva_1[5]), m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_o_expo_mux_11_nl), FpAdd_6U_10U_1_mux_3_itm);
  assign FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_nl = ~(m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_1_mux_3_itm));
  assign FpAdd_6U_10U_1_o_expo_and_7_nl = m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_1_mux_3_itm;
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3,
      (FpAdd_6U_10U_1_o_expo_1_sva_1[3:0]), (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_nl) , (FpAdd_6U_10U_1_o_expo_and_7_nl)
      , (~ FpAdd_6U_10U_1_mux_3_itm)});
  assign FpAdd_6U_10U_1_o_expo_mux_13_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_1_o_expo_1_sva_1[4]), m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_o_expo_mux_13_nl), FpAdd_6U_10U_1_mux_3_itm);
  assign nl_m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_1_mux_3_itm);
  assign FpMantRNE_23U_11U_1_else_carry_1_sva = (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_1_o_expo_1_sva_1 = ({reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_1_sva_1 = nl_FpAdd_6U_10U_1_o_expo_1_sva_1[5:0];
  assign FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row1_1_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_9);
  assign FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_1_int_mant_p1_1_sva_1[22:0]),
      (FpAdd_6U_10U_1_int_mant_p1_1_sva[22:0]), reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_1_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_1_sva, reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign nl_m_row1_1_FpNormalize_6U_23U_1_else_acc_nl = ({reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_36)})
      + 6'b1;
  assign m_row1_1_FpNormalize_6U_23U_1_else_acc_nl = nl_m_row1_1_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row1_1_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_9);
  assign nl_FpAdd_6U_10U_1_o_expo_1_sva_4 = ({FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_1_sva_4 = nl_FpAdd_6U_10U_1_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl = FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm
      | (~ m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl), m_row1_1_FpMantRNE_23U_11U_1_else_and_tmp);
  assign nl_m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl = nl_m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl[5:0];
  assign m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm = ~(m_row1_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1[23])));
  assign nl_m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_1_sva);
  assign m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl = nl_m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_4_itm = MUX_v_10_2_2((m_row1_1_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_2_sva = nl_FpAdd_6U_10U_1_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_1_a_int_mant_p1_2_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_2_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1[23:0];
  assign FpAdd_6U_10U_1_o_expo_mux_17_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_1_o_expo_2_sva_1[5]), m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_o_expo_mux_17_nl), FpAdd_6U_10U_1_mux_20_itm);
  assign FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_1_nl = ~(m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_1_mux_20_itm));
  assign FpAdd_6U_10U_1_o_expo_and_5_nl = m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_1_mux_20_itm;
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3,
      (FpAdd_6U_10U_1_o_expo_2_sva_1[3:0]), (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_1_nl) , (FpAdd_6U_10U_1_o_expo_and_5_nl)
      , (~ FpAdd_6U_10U_1_mux_20_itm)});
  assign FpAdd_6U_10U_1_o_expo_mux_19_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_1_o_expo_2_sva_1[4]), m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_o_expo_mux_19_nl), FpAdd_6U_10U_1_mux_20_itm);
  assign nl_m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_1_mux_20_itm);
  assign FpMantRNE_23U_11U_1_else_carry_2_sva = (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_1_o_expo_2_sva_1 = ({reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_2_sva_1 = nl_FpAdd_6U_10U_1_o_expo_2_sva_1[5:0];
  assign FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row1_2_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_11);
  assign FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_1_int_mant_p1_2_sva_1[22:0]),
      (FpAdd_6U_10U_1_int_mant_p1_2_sva[22:0]), reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_2_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_2_sva, reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign nl_m_row1_2_FpNormalize_6U_23U_1_else_acc_nl = ({reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_37)})
      + 6'b1;
  assign m_row1_2_FpNormalize_6U_23U_1_else_acc_nl = nl_m_row1_2_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row1_2_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_11);
  assign nl_FpAdd_6U_10U_1_o_expo_2_sva_4 = ({FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_2_sva_4 = nl_FpAdd_6U_10U_1_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl = FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm
      | (~ m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl), m_row1_2_FpMantRNE_23U_11U_1_else_and_tmp);
  assign nl_m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl = nl_m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl[5:0];
  assign m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm = ~(m_row1_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1[23])));
  assign nl_m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_2_sva);
  assign m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl = nl_m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_5_itm = MUX_v_10_2_2((m_row1_2_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_3_sva = nl_FpAdd_6U_10U_1_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_1_a_int_mant_p1_3_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_3_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1[23:0];
  assign FpAdd_6U_10U_1_o_expo_mux_23_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_1_o_expo_3_sva_1[5]), m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_o_expo_mux_23_nl), FpAdd_6U_10U_1_mux_37_itm);
  assign FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_2_nl = ~(m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_1_mux_37_itm));
  assign FpAdd_6U_10U_1_o_expo_and_3_nl = m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_1_mux_37_itm;
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3,
      (FpAdd_6U_10U_1_o_expo_3_sva_1[3:0]), (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_2_nl) , (FpAdd_6U_10U_1_o_expo_and_3_nl)
      , (~ FpAdd_6U_10U_1_mux_37_itm)});
  assign FpAdd_6U_10U_1_o_expo_mux_25_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_1_o_expo_3_sva_1[4]), m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_o_expo_mux_25_nl), FpAdd_6U_10U_1_mux_37_itm);
  assign nl_m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_1_mux_37_itm);
  assign FpMantRNE_23U_11U_1_else_carry_3_sva = (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_1_o_expo_3_sva_1 = ({reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_3_sva_1 = nl_FpAdd_6U_10U_1_o_expo_3_sva_1[5:0];
  assign FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row1_3_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_13);
  assign FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_1_int_mant_p1_3_sva_1[22:0]),
      (FpAdd_6U_10U_1_int_mant_p1_3_sva[22:0]), reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_3_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_3_sva, reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign nl_m_row1_3_FpNormalize_6U_23U_1_else_acc_nl = ({reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_38)})
      + 6'b1;
  assign m_row1_3_FpNormalize_6U_23U_1_else_acc_nl = nl_m_row1_3_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row1_3_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_13);
  assign nl_FpAdd_6U_10U_1_o_expo_3_sva_4 = ({FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_3_sva_4 = nl_FpAdd_6U_10U_1_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl = FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm
      | (~ m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl), m_row1_3_FpMantRNE_23U_11U_1_else_and_tmp);
  assign nl_m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl = nl_m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl[5:0];
  assign m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm = ~(m_row1_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1[23])));
  assign nl_m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_3_sva);
  assign m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl = nl_m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_6_itm = MUX_v_10_2_2((m_row1_3_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_sva = nl_FpAdd_6U_10U_1_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_sva_2,
      FpAdd_6U_10U_1_a_int_mant_p1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_sva_2,
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_sva_1[23:0];
  assign FpAdd_6U_10U_1_o_expo_mux_29_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_1_o_expo_sva_1[5]), m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_o_expo_mux_29_nl), FpAdd_6U_10U_1_mux_73_itm);
  assign FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_3_nl = ~(m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_1_mux_73_itm));
  assign FpAdd_6U_10U_1_o_expo_and_1_nl = m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_1_mux_73_itm;
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3,
      (FpAdd_6U_10U_1_o_expo_sva_1[3:0]), (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_1_o_expo_FpAdd_6U_10U_1_o_expo_nor_3_nl) , (FpAdd_6U_10U_1_o_expo_and_1_nl)
      , (~ FpAdd_6U_10U_1_mux_73_itm)});
  assign FpAdd_6U_10U_1_o_expo_mux_31_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_1_o_expo_sva_1[4]), m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_o_expo_mux_31_nl), FpAdd_6U_10U_1_mux_73_itm);
  assign nl_FpAdd_6U_10U_1_o_expo_sva_1 = ({reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_sva_1 = nl_FpAdd_6U_10U_1_o_expo_sva_1[5:0];
  assign nl_m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row1_4_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_15);
  assign FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_1_int_mant_p1_sva_1[22:0]),
      (FpAdd_6U_10U_1_int_mant_p1_sva[22:0]), reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_sva, reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign nl_m_row1_4_FpNormalize_6U_23U_1_else_acc_nl = ({reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_39)})
      + 6'b1;
  assign m_row1_4_FpNormalize_6U_23U_1_else_acc_nl = nl_m_row1_4_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row1_4_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_15);
  assign nl_m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl = nl_m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl[5:0];
  assign m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_2_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_2_int_mant_p1_1_sva = nl_FpAdd_6U_10U_2_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_2_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_2_a_int_mant_p1_1_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_2_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_2_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_2_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_2_int_mant_p1_1_sva_1 = nl_FpAdd_6U_10U_2_int_mant_p1_1_sva_1[23:0];
  assign FpAdd_6U_10U_2_o_expo_mux_11_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_2_o_expo_1_sva_1[5]), m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_2_o_expo_mux_11_nl), FpAdd_6U_10U_2_mux_3_itm);
  assign FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_nl = ~(m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_2_mux_3_itm));
  assign FpAdd_6U_10U_2_o_expo_and_7_nl = m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_2_mux_3_itm;
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3,
      (FpAdd_6U_10U_2_o_expo_1_sva_1[3:0]), (FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_nl) , (FpAdd_6U_10U_2_o_expo_and_7_nl)
      , (~ FpAdd_6U_10U_2_mux_3_itm)});
  assign FpAdd_6U_10U_2_o_expo_mux_13_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_2_o_expo_1_sva_1[4]), m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_2_o_expo_mux_13_nl), FpAdd_6U_10U_2_mux_3_itm);
  assign nl_m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl = nl_m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl[5:0];
  assign m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_2_mux_3_itm);
  assign FpMantRNE_23U_11U_2_else_carry_1_sva = (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_2_o_expo_1_sva_1 = ({reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_1_sva_1 = nl_FpAdd_6U_10U_2_o_expo_1_sva_1[5:0];
  assign FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row2_1_FpNormalize_6U_23U_2_else_lshift_itm, FpNormalize_6U_23U_2_oelse_not_9);
  assign FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_2_int_mant_p1_1_sva_1[22:0]),
      (FpAdd_6U_10U_2_int_mant_p1_1_sva[22:0]), reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_2_int_mant_p1_1_sva_1,
      FpAdd_6U_10U_2_int_mant_p1_1_sva, reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign nl_m_row2_1_FpNormalize_6U_23U_2_else_acc_nl = ({reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_40)})
      + 6'b1;
  assign m_row2_1_FpNormalize_6U_23U_2_else_acc_nl = nl_m_row2_1_FpNormalize_6U_23U_2_else_acc_nl[5:0];
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row2_1_FpNormalize_6U_23U_2_else_acc_nl),
      FpNormalize_6U_23U_2_oelse_not_9);
  assign nl_FpAdd_6U_10U_2_o_expo_1_sva_4 = ({FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_1_sva_4 = nl_FpAdd_6U_10U_2_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_nl = FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm
      | (~ m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_nl), m_row2_1_FpMantRNE_23U_11U_2_else_and_tmp);
  assign nl_m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl = nl_m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl[5:0];
  assign m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm = ~(m_row2_1_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1[23])));
  assign nl_m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl = (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_2_else_carry_1_sva);
  assign m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl = nl_m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl[9:0];
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_4_itm = MUX_v_10_2_2((m_row2_1_FpMantRNE_23U_11U_2_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_2_int_mant_p1_2_sva = nl_FpAdd_6U_10U_2_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_2_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_2_a_int_mant_p1_2_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_2_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_2_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_2_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_2_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_2_int_mant_p1_2_sva_1 = nl_FpAdd_6U_10U_2_int_mant_p1_2_sva_1[23:0];
  assign FpAdd_6U_10U_2_o_expo_mux_17_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_2_o_expo_2_sva_1[5]), m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_2_o_expo_mux_17_nl), FpAdd_6U_10U_2_mux_20_itm);
  assign FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_1_nl = ~(m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_2_mux_20_itm));
  assign FpAdd_6U_10U_2_o_expo_and_5_nl = m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_2_mux_20_itm;
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3,
      (FpAdd_6U_10U_2_o_expo_2_sva_1[3:0]), (FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_1_nl) , (FpAdd_6U_10U_2_o_expo_and_5_nl)
      , (~ FpAdd_6U_10U_2_mux_20_itm)});
  assign FpAdd_6U_10U_2_o_expo_mux_19_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_2_o_expo_2_sva_1[4]), m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_2_o_expo_mux_19_nl), FpAdd_6U_10U_2_mux_20_itm);
  assign nl_m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl = nl_m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl[5:0];
  assign m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_2_mux_20_itm);
  assign FpMantRNE_23U_11U_2_else_carry_2_sva = (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_2_o_expo_2_sva_1 = ({reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_2_sva_1 = nl_FpAdd_6U_10U_2_o_expo_2_sva_1[5:0];
  assign FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row2_2_FpNormalize_6U_23U_2_else_lshift_itm, FpNormalize_6U_23U_2_oelse_not_11);
  assign FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_2_int_mant_p1_2_sva_1[22:0]),
      (FpAdd_6U_10U_2_int_mant_p1_2_sva[22:0]), reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_2_int_mant_p1_2_sva_1,
      FpAdd_6U_10U_2_int_mant_p1_2_sva, reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign nl_m_row2_2_FpNormalize_6U_23U_2_else_acc_nl = ({reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_41)})
      + 6'b1;
  assign m_row2_2_FpNormalize_6U_23U_2_else_acc_nl = nl_m_row2_2_FpNormalize_6U_23U_2_else_acc_nl[5:0];
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row2_2_FpNormalize_6U_23U_2_else_acc_nl),
      FpNormalize_6U_23U_2_oelse_not_11);
  assign nl_FpAdd_6U_10U_2_o_expo_2_sva_4 = ({FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_2_sva_4 = nl_FpAdd_6U_10U_2_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_1_nl = FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm
      | (~ m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_1_nl), m_row2_2_FpMantRNE_23U_11U_2_else_and_tmp);
  assign nl_m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl = nl_m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl[5:0];
  assign m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm = ~(m_row2_2_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1[23])));
  assign nl_m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl = (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_2_else_carry_2_sva);
  assign m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl = nl_m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl[9:0];
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_5_itm = MUX_v_10_2_2((m_row2_2_FpMantRNE_23U_11U_2_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_2_int_mant_p1_3_sva = nl_FpAdd_6U_10U_2_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_2_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_2_a_int_mant_p1_3_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_2_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_2_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_3_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_2_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_2_int_mant_p1_3_sva_1 = nl_FpAdd_6U_10U_2_int_mant_p1_3_sva_1[23:0];
  assign FpAdd_6U_10U_2_o_expo_mux_23_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_2_o_expo_3_sva_1[5]), m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_2_o_expo_mux_23_nl), FpAdd_6U_10U_2_mux_37_itm);
  assign FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_2_nl = ~(m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_2_mux_37_itm));
  assign FpAdd_6U_10U_2_o_expo_and_3_nl = m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_2_mux_37_itm;
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3,
      (FpAdd_6U_10U_2_o_expo_3_sva_1[3:0]), (FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_2_nl) , (FpAdd_6U_10U_2_o_expo_and_3_nl)
      , (~ FpAdd_6U_10U_2_mux_37_itm)});
  assign FpAdd_6U_10U_2_o_expo_mux_25_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_2_o_expo_3_sva_1[4]), m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_2_o_expo_mux_25_nl), FpAdd_6U_10U_2_mux_37_itm);
  assign nl_m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl = nl_m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl[5:0];
  assign m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_2_mux_37_itm);
  assign FpMantRNE_23U_11U_2_else_carry_3_sva = (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_2_o_expo_3_sva_1 = ({reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_3_sva_1 = nl_FpAdd_6U_10U_2_o_expo_3_sva_1[5:0];
  assign FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row2_3_FpNormalize_6U_23U_2_else_lshift_itm, FpNormalize_6U_23U_2_oelse_not_13);
  assign FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_2_int_mant_p1_3_sva_1[22:0]),
      (FpAdd_6U_10U_2_int_mant_p1_3_sva[22:0]), reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_2_int_mant_p1_3_sva_1,
      FpAdd_6U_10U_2_int_mant_p1_3_sva, reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign nl_m_row2_3_FpNormalize_6U_23U_2_else_acc_nl = ({reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_42)})
      + 6'b1;
  assign m_row2_3_FpNormalize_6U_23U_2_else_acc_nl = nl_m_row2_3_FpNormalize_6U_23U_2_else_acc_nl[5:0];
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row2_3_FpNormalize_6U_23U_2_else_acc_nl),
      FpNormalize_6U_23U_2_oelse_not_13);
  assign nl_FpAdd_6U_10U_2_o_expo_3_sva_4 = ({FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_3_sva_4 = nl_FpAdd_6U_10U_2_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_2_nl = FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm
      | (~ m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_2_nl), m_row2_3_FpMantRNE_23U_11U_2_else_and_tmp);
  assign nl_m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl = nl_m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl[5:0];
  assign m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm = ~(m_row2_3_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1[23])));
  assign nl_m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl = (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_2_else_carry_3_sva);
  assign m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl = nl_m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl[9:0];
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_6_itm = MUX_v_10_2_2((m_row2_3_FpMantRNE_23U_11U_2_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_2_int_mant_p1_sva = nl_FpAdd_6U_10U_2_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_2_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_sva_2,
      FpAdd_6U_10U_2_a_int_mant_p1_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_6U_10U_2_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_sva_2,
      FpAdd_6U_10U_2_b_int_mant_p1_sva_2, FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_2_int_mant_p1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_2_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_2_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_2_int_mant_p1_sva_1 = nl_FpAdd_6U_10U_2_int_mant_p1_sva_1[23:0];
  assign FpAdd_6U_10U_2_o_expo_mux_29_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_2_o_expo_sva_1[5]), m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_2_o_expo_mux_29_nl), FpAdd_6U_10U_2_mux_73_itm);
  assign FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_3_nl = ~(m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_2_mux_73_itm));
  assign FpAdd_6U_10U_2_o_expo_and_1_nl = m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_2_mux_73_itm;
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3,
      (FpAdd_6U_10U_2_o_expo_sva_1[3:0]), (FpAdd_6U_10U_2_o_expo_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_2_o_expo_FpAdd_6U_10U_2_o_expo_nor_3_nl) , (FpAdd_6U_10U_2_o_expo_and_1_nl)
      , (~ FpAdd_6U_10U_2_mux_73_itm)});
  assign FpAdd_6U_10U_2_o_expo_mux_31_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_2_o_expo_sva_1[4]), m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_2_o_expo_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_2_o_expo_mux_31_nl), FpAdd_6U_10U_2_mux_73_itm);
  assign nl_FpAdd_6U_10U_2_o_expo_sva_1 = ({reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_sva_1 = nl_FpAdd_6U_10U_2_o_expo_sva_1[5:0];
  assign nl_m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl = nl_m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl[5:0];
  assign m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row2_4_FpNormalize_6U_23U_2_else_lshift_itm, FpNormalize_6U_23U_2_oelse_not_15);
  assign FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_2_int_mant_p1_sva_1[22:0]),
      (FpAdd_6U_10U_2_int_mant_p1_sva[22:0]), reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_2_int_mant_p1_sva_1,
      FpAdd_6U_10U_2_int_mant_p1_sva, reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign nl_m_row2_4_FpNormalize_6U_23U_2_else_acc_nl = ({reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_43)})
      + 6'b1;
  assign m_row2_4_FpNormalize_6U_23U_2_else_acc_nl = nl_m_row2_4_FpNormalize_6U_23U_2_else_acc_nl[5:0];
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row2_4_FpNormalize_6U_23U_2_else_acc_nl),
      FpNormalize_6U_23U_2_oelse_not_15);
  assign nl_m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl = nl_m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl[5:0];
  assign m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_3_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_3_int_mant_p1_1_sva = nl_FpAdd_6U_10U_3_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_3_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_3_a_int_mant_p1_1_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_4);
  assign FpAdd_6U_10U_3_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_3_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_3_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_3_int_mant_p1_1_sva_1 = nl_FpAdd_6U_10U_3_int_mant_p1_1_sva_1[23:0];
  assign FpAdd_6U_10U_3_o_expo_mux_11_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_3_o_expo_1_sva_1[5]), m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_3_o_expo_mux_11_nl), FpAdd_6U_10U_3_mux_3_itm);
  assign FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_nl = ~(m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_3_mux_3_itm));
  assign FpAdd_6U_10U_3_o_expo_and_7_nl = m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_3_mux_3_itm;
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3,
      (FpAdd_6U_10U_3_o_expo_1_sva_1[3:0]), (FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_nl) , (FpAdd_6U_10U_3_o_expo_and_7_nl)
      , (~ FpAdd_6U_10U_3_mux_3_itm)});
  assign FpAdd_6U_10U_3_o_expo_mux_13_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_3_o_expo_1_sva_1[4]), m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_3_o_expo_mux_13_nl), FpAdd_6U_10U_3_mux_3_itm);
  assign nl_m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl = nl_m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl[5:0];
  assign m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_3_mux_3_itm);
  assign FpMantRNE_23U_11U_3_else_carry_1_sva = (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_3_o_expo_1_sva_1 = ({reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_1_sva_1 = nl_FpAdd_6U_10U_3_o_expo_1_sva_1[5:0];
  assign FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row3_1_FpNormalize_6U_23U_3_else_lshift_itm, FpNormalize_6U_23U_3_oelse_not_9);
  assign FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_3_int_mant_p1_1_sva_1[22:0]),
      (FpAdd_6U_10U_3_int_mant_p1_1_sva[22:0]), reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_3_int_mant_p1_1_sva_1,
      FpAdd_6U_10U_3_int_mant_p1_1_sva, reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign nl_m_row3_1_FpNormalize_6U_23U_3_else_acc_nl = ({reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_44)})
      + 6'b1;
  assign m_row3_1_FpNormalize_6U_23U_3_else_acc_nl = nl_m_row3_1_FpNormalize_6U_23U_3_else_acc_nl[5:0];
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row3_1_FpNormalize_6U_23U_3_else_acc_nl),
      FpNormalize_6U_23U_3_oelse_not_9);
  assign nl_FpAdd_6U_10U_3_o_expo_1_sva_4 = ({FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_1_sva_4 = nl_FpAdd_6U_10U_3_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_nl = FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm
      | (~ m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_nl), m_row3_1_FpMantRNE_23U_11U_3_else_and_tmp);
  assign nl_m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl = nl_m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl[5:0];
  assign m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm = ~(m_row3_1_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1[23])));
  assign nl_m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl = (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_3_else_carry_1_sva);
  assign m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl = nl_m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl[9:0];
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_4_itm = MUX_v_10_2_2((m_row3_1_FpMantRNE_23U_11U_3_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_3_int_mant_p1_2_sva = nl_FpAdd_6U_10U_3_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_3_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_3_a_int_mant_p1_2_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_4);
  assign FpAdd_6U_10U_3_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_3_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_2_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_3_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_3_int_mant_p1_2_sva_1 = nl_FpAdd_6U_10U_3_int_mant_p1_2_sva_1[23:0];
  assign FpAdd_6U_10U_3_o_expo_mux_17_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_3_o_expo_2_sva_1[5]), m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_3_o_expo_mux_17_nl), FpAdd_6U_10U_3_mux_20_itm);
  assign FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_1_nl = ~(m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_3_mux_20_itm));
  assign FpAdd_6U_10U_3_o_expo_and_5_nl = m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_3_mux_20_itm;
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3,
      (FpAdd_6U_10U_3_o_expo_2_sva_1[3:0]), (FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_1_nl) , (FpAdd_6U_10U_3_o_expo_and_5_nl)
      , (~ FpAdd_6U_10U_3_mux_20_itm)});
  assign FpAdd_6U_10U_3_o_expo_mux_19_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_3_o_expo_2_sva_1[4]), m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_3_o_expo_mux_19_nl), FpAdd_6U_10U_3_mux_20_itm);
  assign nl_m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl = nl_m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl[5:0];
  assign m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_3_mux_20_itm);
  assign FpMantRNE_23U_11U_3_else_carry_2_sva = (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_3_o_expo_2_sva_1 = ({reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_2_sva_1 = nl_FpAdd_6U_10U_3_o_expo_2_sva_1[5:0];
  assign FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row3_2_FpNormalize_6U_23U_3_else_lshift_itm, FpNormalize_6U_23U_3_oelse_not_11);
  assign FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_3_int_mant_p1_2_sva_1[22:0]),
      (FpAdd_6U_10U_3_int_mant_p1_2_sva[22:0]), reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_3_int_mant_p1_2_sva_1,
      FpAdd_6U_10U_3_int_mant_p1_2_sva, reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign nl_m_row3_2_FpNormalize_6U_23U_3_else_acc_nl = ({reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_45)})
      + 6'b1;
  assign m_row3_2_FpNormalize_6U_23U_3_else_acc_nl = nl_m_row3_2_FpNormalize_6U_23U_3_else_acc_nl[5:0];
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row3_2_FpNormalize_6U_23U_3_else_acc_nl),
      FpNormalize_6U_23U_3_oelse_not_11);
  assign nl_FpAdd_6U_10U_3_o_expo_2_sva_4 = ({FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_2_sva_4 = nl_FpAdd_6U_10U_3_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_1_nl = FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm
      | (~ m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_1_nl), m_row3_2_FpMantRNE_23U_11U_3_else_and_tmp);
  assign nl_m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl = nl_m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl[5:0];
  assign m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm = ~(m_row3_2_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1[23])));
  assign nl_m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl = (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_3_else_carry_2_sva);
  assign m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl = nl_m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl[9:0];
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_5_itm = MUX_v_10_2_2((m_row3_2_FpMantRNE_23U_11U_3_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_3_int_mant_p1_3_sva = nl_FpAdd_6U_10U_3_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_3_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_3_a_int_mant_p1_3_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_4);
  assign FpAdd_6U_10U_3_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_3_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_3_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_3_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_3_int_mant_p1_3_sva_1 = nl_FpAdd_6U_10U_3_int_mant_p1_3_sva_1[23:0];
  assign FpAdd_6U_10U_3_o_expo_mux_23_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_3_o_expo_3_sva_1[5]), m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_3_o_expo_mux_23_nl), FpAdd_6U_10U_3_mux_37_itm);
  assign FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_2_nl = ~(m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_3_mux_37_itm));
  assign FpAdd_6U_10U_3_o_expo_and_3_nl = m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_3_mux_37_itm;
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3,
      (FpAdd_6U_10U_3_o_expo_3_sva_1[3:0]), (FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_2_nl) , (FpAdd_6U_10U_3_o_expo_and_3_nl)
      , (~ FpAdd_6U_10U_3_mux_37_itm)});
  assign FpAdd_6U_10U_3_o_expo_mux_25_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_3_o_expo_3_sva_1[4]), m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_3_o_expo_mux_25_nl), FpAdd_6U_10U_3_mux_37_itm);
  assign nl_m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl = nl_m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl[5:0];
  assign m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_3_mux_37_itm);
  assign FpMantRNE_23U_11U_3_else_carry_3_sva = (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign nl_FpAdd_6U_10U_3_o_expo_3_sva_1 = ({reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_3_sva_1 = nl_FpAdd_6U_10U_3_o_expo_3_sva_1[5:0];
  assign FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row3_3_FpNormalize_6U_23U_3_else_lshift_itm, FpNormalize_6U_23U_3_oelse_not_13);
  assign FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_3_int_mant_p1_3_sva_1[22:0]),
      (FpAdd_6U_10U_3_int_mant_p1_3_sva[22:0]), reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_3_int_mant_p1_3_sva_1,
      FpAdd_6U_10U_3_int_mant_p1_3_sva, reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign nl_m_row3_3_FpNormalize_6U_23U_3_else_acc_nl = ({reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_46)})
      + 6'b1;
  assign m_row3_3_FpNormalize_6U_23U_3_else_acc_nl = nl_m_row3_3_FpNormalize_6U_23U_3_else_acc_nl[5:0];
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row3_3_FpNormalize_6U_23U_3_else_acc_nl),
      FpNormalize_6U_23U_3_oelse_not_13);
  assign nl_FpAdd_6U_10U_3_o_expo_3_sva_4 = ({FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_3_sva_4 = nl_FpAdd_6U_10U_3_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_2_nl = FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm
      | (~ m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_2_nl), m_row3_3_FpMantRNE_23U_11U_3_else_and_tmp);
  assign nl_m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl = nl_m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl[5:0];
  assign m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm = ~(m_row3_3_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1[23])));
  assign nl_m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl = (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_3_else_carry_3_sva);
  assign m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl = nl_m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl[9:0];
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_6_itm = MUX_v_10_2_2((m_row3_3_FpMantRNE_23U_11U_3_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_3_int_mant_p1_sva = nl_FpAdd_6U_10U_3_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_3_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_sva_2,
      FpAdd_6U_10U_3_a_int_mant_p1_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_4);
  assign FpAdd_6U_10U_3_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_sva_2,
      FpAdd_6U_10U_3_b_int_mant_p1_sva_2, FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_4);
  assign nl_FpAdd_6U_10U_3_int_mant_p1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_3_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_3_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_3_int_mant_p1_sva_1 = nl_FpAdd_6U_10U_3_int_mant_p1_sva_1[23:0];
  assign FpAdd_6U_10U_3_o_expo_mux_29_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp,
      (FpAdd_6U_10U_3_o_expo_sva_1[5]), m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_5_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_3_o_expo_mux_29_nl), FpAdd_6U_10U_3_mux_69_itm);
  assign FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_3_nl = ~(m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ FpAdd_6U_10U_3_mux_69_itm));
  assign FpAdd_6U_10U_3_o_expo_and_1_nl = m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      & FpAdd_6U_10U_3_mux_69_itm;
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_3_0_mx0 = MUX1HOT_v_4_3_2(FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3,
      (FpAdd_6U_10U_3_o_expo_sva_1[3:0]), (FpAdd_6U_10U_3_o_expo_lpi_1_dfm_1[3:0]),
      {(FpAdd_6U_10U_3_o_expo_FpAdd_6U_10U_3_o_expo_nor_3_nl) , (FpAdd_6U_10U_3_o_expo_and_1_nl)
      , (~ FpAdd_6U_10U_3_mux_69_itm)});
  assign FpAdd_6U_10U_3_o_expo_mux_31_nl = MUX_s_1_2_2(reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1,
      (FpAdd_6U_10U_3_o_expo_sva_1[4]), m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_4_mx0 = MUX_s_1_2_2((FpAdd_6U_10U_3_o_expo_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_3_o_expo_mux_31_nl), FpAdd_6U_10U_3_mux_69_itm);
  assign nl_FpAdd_6U_10U_3_o_expo_sva_1 = ({reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_sva_1 = nl_FpAdd_6U_10U_3_o_expo_sva_1[5:0];
  assign nl_m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1 , (FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3[3:1])})
      + 6'b1;
  assign m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl = nl_m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl[5:0];
  assign m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      m_row3_4_FpNormalize_6U_23U_3_else_lshift_itm, FpNormalize_6U_23U_3_oelse_not_15);
  assign FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx0_tmp_22_0 = MUX_v_23_2_2((FpAdd_6U_10U_3_int_mant_p1_sva_1[22:0]),
      (FpAdd_6U_10U_3_int_mant_p1_sva[22:0]), reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1 = MUX_v_24_2_2(FpAdd_6U_10U_3_int_mant_p1_sva_1,
      FpAdd_6U_10U_3_int_mant_p1_sva, reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign nl_m_row3_4_FpNormalize_6U_23U_3_else_acc_nl = ({reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1 , FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_47)})
      + 6'b1;
  assign m_row3_4_FpNormalize_6U_23U_3_else_acc_nl = nl_m_row3_4_FpNormalize_6U_23U_3_else_acc_nl[5:0];
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (m_row3_4_FpNormalize_6U_23U_3_else_acc_nl),
      FpNormalize_6U_23U_3_oelse_not_15);
  assign nl_m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_4_mx0 , (FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_3_0_mx0[3:1])})
      + 6'b1;
  assign m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl = nl_m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl[5:0];
  assign m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse = IsNaN_6U_10U_7_land_3_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_6_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse);
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_13_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_3_o_expo_3_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse , FpAdd_6U_10U_3_and_24_ssc
      , FpAdd_6U_10U_3_and_17_ssc});
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_5 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_13_nl)
      | FpAdd_6U_10U_3_and_25_ssc;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_2_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_3_o_expo_3_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse , FpAdd_6U_10U_3_and_24_ssc
      , FpAdd_6U_10U_3_and_17_ssc});
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_4 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_2_nl)
      | FpAdd_6U_10U_3_and_25_ssc;
  assign FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_7,
      FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_3_o_expo_3_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse , FpAdd_6U_10U_3_and_24_ssc
      , FpAdd_6U_10U_3_and_17_ssc , FpAdd_6U_10U_3_and_25_ssc});
  assign FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_6_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_7, or_1963_cse);
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_13_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_2_o_expo_3_sva_4[5]),
      {or_1963_cse , FpAdd_6U_10U_2_and_24_ssc , FpAdd_6U_10U_2_and_17_ssc});
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_5 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_13_nl)
      | FpAdd_6U_10U_2_and_25_ssc;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_2_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_2_o_expo_3_sva_4[4]),
      {or_1963_cse , FpAdd_6U_10U_2_and_24_ssc , FpAdd_6U_10U_2_and_17_ssc});
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_4 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_2_nl)
      | FpAdd_6U_10U_2_and_25_ssc;
  assign FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_7,
      FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_2_o_expo_3_sva_4[3:0]),
      4'b1110, {or_1963_cse , FpAdd_6U_10U_2_and_24_ssc , FpAdd_6U_10U_2_and_17_ssc
      , FpAdd_6U_10U_2_and_25_ssc});
  assign FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_6_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7, or_1960_cse);
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_13_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_1_o_expo_3_sva_4[5]),
      {or_1960_cse , FpAdd_6U_10U_1_and_24_ssc , FpAdd_6U_10U_1_and_17_ssc});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_13_nl)
      | FpAdd_6U_10U_1_and_25_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_1_o_expo_3_sva_4[4]),
      {or_1960_cse , FpAdd_6U_10U_1_and_24_ssc , FpAdd_6U_10U_1_and_17_ssc});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl)
      | FpAdd_6U_10U_1_and_25_ssc;
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_7,
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_1_o_expo_3_sva_4[3:0]),
      4'b1110, {or_1960_cse , FpAdd_6U_10U_1_and_24_ssc , FpAdd_6U_10U_1_and_17_ssc
      , FpAdd_6U_10U_1_and_25_ssc});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse = IsNaN_6U_10U_1_land_3_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_FpAdd_6U_10U_or_6_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse);
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_o_expo_3_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse , FpAdd_6U_10U_and_24_ssc
      , FpAdd_6U_10U_and_17_ssc});
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl)
      | FpAdd_6U_10U_and_25_ssc;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_2_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_o_expo_3_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse , FpAdd_6U_10U_and_24_ssc
      , FpAdd_6U_10U_and_17_ssc});
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_4 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_2_nl)
      | FpAdd_6U_10U_and_25_ssc;
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_7,
      FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_o_expo_3_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse , FpAdd_6U_10U_and_24_ssc
      , FpAdd_6U_10U_and_17_ssc , FpAdd_6U_10U_and_25_ssc});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse = IsNaN_6U_10U_7_land_2_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse);
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_11_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_3_o_expo_2_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse , FpAdd_6U_10U_3_and_22_ssc
      , FpAdd_6U_10U_3_and_15_ssc});
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_5 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_11_nl)
      | FpAdd_6U_10U_3_and_23_ssc;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_1_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_3_o_expo_2_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse , FpAdd_6U_10U_3_and_22_ssc
      , FpAdd_6U_10U_3_and_15_ssc});
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_4 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_1_nl)
      | FpAdd_6U_10U_3_and_23_ssc;
  assign FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_7,
      FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_3_o_expo_2_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse , FpAdd_6U_10U_3_and_22_ssc
      , FpAdd_6U_10U_3_and_15_ssc , FpAdd_6U_10U_3_and_23_ssc});
  assign FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_7, or_1962_cse);
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_11_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_2_o_expo_2_sva_4[5]),
      {or_1962_cse , FpAdd_6U_10U_2_and_22_ssc , FpAdd_6U_10U_2_and_15_ssc});
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_5 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_11_nl)
      | FpAdd_6U_10U_2_and_23_ssc;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_1_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_2_o_expo_2_sva_4[4]),
      {or_1962_cse , FpAdd_6U_10U_2_and_22_ssc , FpAdd_6U_10U_2_and_15_ssc});
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_4 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_1_nl)
      | FpAdd_6U_10U_2_and_23_ssc;
  assign FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_7,
      FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_2_o_expo_2_sva_4[3:0]),
      4'b1110, {or_1962_cse , FpAdd_6U_10U_2_and_22_ssc , FpAdd_6U_10U_2_and_15_ssc
      , FpAdd_6U_10U_2_and_23_ssc});
  assign IsNaN_6U_10U_10_nor_1_tmp = ~((FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000));
  assign IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp = ~(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5
      & FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4 & (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0==4'b1111));
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_1_o_expo_2_sva_4[5]),
      {or_1959_cse , FpAdd_6U_10U_1_and_22_ssc , FpAdd_6U_10U_1_and_15_ssc});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl)
      | FpAdd_6U_10U_1_and_23_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_1_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_1_o_expo_2_sva_4[4]),
      {or_1959_cse , FpAdd_6U_10U_1_and_22_ssc , FpAdd_6U_10U_1_and_15_ssc});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_1_nl)
      | FpAdd_6U_10U_1_and_23_ssc;
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_7,
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_1_o_expo_2_sva_4[3:0]),
      4'b1110, {or_1959_cse , FpAdd_6U_10U_1_and_22_ssc , FpAdd_6U_10U_1_and_15_ssc
      , FpAdd_6U_10U_1_and_23_ssc});
  assign FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_7, or_1959_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse = IsNaN_6U_10U_1_land_2_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_FpAdd_6U_10U_or_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse);
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_11_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_o_expo_2_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse , FpAdd_6U_10U_and_22_ssc
      , FpAdd_6U_10U_and_15_ssc});
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_11_nl)
      | FpAdd_6U_10U_and_23_ssc;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_1_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_o_expo_2_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse , FpAdd_6U_10U_and_22_ssc
      , FpAdd_6U_10U_and_15_ssc});
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_4 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_1_nl)
      | FpAdd_6U_10U_and_23_ssc;
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_7,
      FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_o_expo_2_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse , FpAdd_6U_10U_and_22_ssc
      , FpAdd_6U_10U_and_15_ssc , FpAdd_6U_10U_and_23_ssc});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse = IsNaN_6U_10U_7_land_1_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_4_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse);
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_9_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_3_o_expo_1_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse , FpAdd_6U_10U_3_and_20_ssc
      , FpAdd_6U_10U_3_and_13_ssc});
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_5 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_9_nl)
      | FpAdd_6U_10U_3_and_21_ssc;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_3_o_expo_1_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse , FpAdd_6U_10U_3_and_20_ssc
      , FpAdd_6U_10U_3_and_13_ssc});
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_4 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_nl)
      | FpAdd_6U_10U_3_and_21_ssc;
  assign FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_7,
      FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_3_o_expo_1_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse , FpAdd_6U_10U_3_and_20_ssc
      , FpAdd_6U_10U_3_and_13_ssc , FpAdd_6U_10U_3_and_21_ssc});
  assign FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_4_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_7, or_1961_cse);
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_9_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_2_o_expo_1_sva_4[5]),
      {or_1961_cse , FpAdd_6U_10U_2_and_20_ssc , FpAdd_6U_10U_2_and_13_ssc});
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_5 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_9_nl)
      | FpAdd_6U_10U_2_and_21_ssc;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_2_o_expo_1_sva_4[4]),
      {or_1961_cse , FpAdd_6U_10U_2_and_20_ssc , FpAdd_6U_10U_2_and_13_ssc});
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_4 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_nl)
      | FpAdd_6U_10U_2_and_21_ssc;
  assign FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_7,
      FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_2_o_expo_1_sva_4[3:0]),
      4'b1110, {or_1961_cse , FpAdd_6U_10U_2_and_20_ssc , FpAdd_6U_10U_2_and_13_ssc
      , FpAdd_6U_10U_2_and_21_ssc});
  assign FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_4_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_7, or_1958_cse);
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_9_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_1_o_expo_1_sva_4[5]),
      {or_1958_cse , FpAdd_6U_10U_1_and_20_ssc , FpAdd_6U_10U_1_and_13_ssc});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_9_nl)
      | FpAdd_6U_10U_1_and_21_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_1_o_expo_1_sva_4[4]),
      {or_1958_cse , FpAdd_6U_10U_1_and_20_ssc , FpAdd_6U_10U_1_and_13_ssc});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_nl)
      | FpAdd_6U_10U_1_and_21_ssc;
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_7,
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_1_o_expo_1_sva_4[3:0]),
      4'b1110, {or_1958_cse , FpAdd_6U_10U_1_and_20_ssc , FpAdd_6U_10U_1_and_13_ssc
      , FpAdd_6U_10U_1_and_21_ssc});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse = IsNaN_6U_10U_1_land_1_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse;
  assign FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_FpAdd_6U_10U_or_4_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_7, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse);
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_9_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_o_expo_1_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse , FpAdd_6U_10U_and_20_ssc
      , FpAdd_6U_10U_and_13_ssc});
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_9_nl)
      | FpAdd_6U_10U_and_21_ssc;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_o_expo_1_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse , FpAdd_6U_10U_and_20_ssc
      , FpAdd_6U_10U_and_13_ssc});
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_4 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_nl)
      | FpAdd_6U_10U_and_21_ssc;
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_7,
      FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_o_expo_1_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse , FpAdd_6U_10U_and_20_ssc
      , FpAdd_6U_10U_and_13_ssc , FpAdd_6U_10U_and_21_ssc});
  assign m_row3_4_FpMantRNE_23U_11U_3_else_and_tmp = FpMantRNE_23U_11U_3_else_carry_sva
      & (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1[23]));
  assign FpMantRNE_23U_11U_3_else_carry_sva = (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_3_mux_69_itm);
  assign FpAdd_6U_10U_3_and_24_ssc = (~(FpAdd_6U_10U_3_and_10_tmp | FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_6_m1c;
  assign FpAdd_6U_10U_3_and_17_ssc = FpAdd_6U_10U_3_and_10_tmp & (~ FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_6_m1c;
  assign FpAdd_6U_10U_3_and_25_ssc = FpAdd_6U_10U_3_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_6_m1c;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_6_m1c = ~(IsNaN_6U_10U_7_land_3_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_3_and_10_tmp = m_row3_3_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1
      & m_row3_3_FpMantRNE_23U_11U_3_else_and_tmp;
  assign m_row3_3_FpMantRNE_23U_11U_3_else_and_tmp = FpMantRNE_23U_11U_3_else_carry_3_sva
      & (FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_3_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_3_and_22_ssc = (~(FpAdd_6U_10U_3_and_9_tmp | FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_5_m1c;
  assign FpAdd_6U_10U_3_and_15_ssc = FpAdd_6U_10U_3_and_9_tmp & (~ FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_5_m1c;
  assign FpAdd_6U_10U_3_and_23_ssc = FpAdd_6U_10U_3_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_5_m1c;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_5_m1c = ~(IsNaN_6U_10U_7_land_2_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_3_and_9_tmp = m_row3_2_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1
      & m_row3_2_FpMantRNE_23U_11U_3_else_and_tmp;
  assign m_row3_2_FpMantRNE_23U_11U_3_else_and_tmp = FpMantRNE_23U_11U_3_else_carry_2_sva
      & (FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_3_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_3_and_20_ssc = (~(FpAdd_6U_10U_3_and_8_tmp | FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_4_m1c;
  assign FpAdd_6U_10U_3_and_13_ssc = FpAdd_6U_10U_3_and_8_tmp & (~ FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_4_m1c;
  assign FpAdd_6U_10U_3_and_21_ssc = FpAdd_6U_10U_3_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_4_m1c;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_4_m1c = ~(IsNaN_6U_10U_7_land_1_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_3_and_8_tmp = m_row3_1_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1
      & m_row3_1_FpMantRNE_23U_11U_3_else_and_tmp;
  assign m_row3_1_FpMantRNE_23U_11U_3_else_and_tmp = FpMantRNE_23U_11U_3_else_carry_1_sva
      & (FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_3_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1[23]));
  assign m_row2_4_FpMantRNE_23U_11U_2_else_and_tmp = FpMantRNE_23U_11U_2_else_carry_sva
      & (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1[23]));
  assign FpMantRNE_23U_11U_2_else_carry_sva = (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_2_mux_73_itm);
  assign FpAdd_6U_10U_2_and_24_ssc = (~(FpAdd_6U_10U_2_and_10_tmp | FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_6_m1c;
  assign FpAdd_6U_10U_2_and_17_ssc = FpAdd_6U_10U_2_and_10_tmp & (~ FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_6_m1c;
  assign FpAdd_6U_10U_2_and_25_ssc = FpAdd_6U_10U_2_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_6_m1c;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_6_m1c = ~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_3
      | IsNaN_6U_10U_4_land_3_lpi_1_dfm_3);
  assign FpAdd_6U_10U_2_and_10_tmp = m_row2_3_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1
      & m_row2_3_FpMantRNE_23U_11U_2_else_and_tmp;
  assign m_row2_3_FpMantRNE_23U_11U_2_else_and_tmp = FpMantRNE_23U_11U_2_else_carry_3_sva
      & (FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_2_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_2_and_22_ssc = (~(FpAdd_6U_10U_2_and_9_tmp | FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_5_m1c;
  assign FpAdd_6U_10U_2_and_15_ssc = FpAdd_6U_10U_2_and_9_tmp & (~ FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_5_m1c;
  assign FpAdd_6U_10U_2_and_23_ssc = FpAdd_6U_10U_2_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_5_m1c;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_5_m1c = ~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_3
      | IsNaN_6U_10U_4_land_2_lpi_1_dfm_3);
  assign FpAdd_6U_10U_2_and_9_tmp = m_row2_2_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1
      & m_row2_2_FpMantRNE_23U_11U_2_else_and_tmp;
  assign m_row2_2_FpMantRNE_23U_11U_2_else_and_tmp = FpMantRNE_23U_11U_2_else_carry_2_sva
      & (FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_2_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_2_and_20_ssc = (~(FpAdd_6U_10U_2_and_8_tmp | FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_4_m1c;
  assign FpAdd_6U_10U_2_and_13_ssc = FpAdd_6U_10U_2_and_8_tmp & (~ FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_4_m1c;
  assign FpAdd_6U_10U_2_and_21_ssc = FpAdd_6U_10U_2_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_4_m1c;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_4_m1c = ~(IsNaN_6U_10U_5_land_1_lpi_1_dfm_3
      | IsNaN_6U_10U_4_land_1_lpi_1_dfm_3);
  assign FpAdd_6U_10U_2_and_8_tmp = m_row2_1_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1
      & m_row2_1_FpMantRNE_23U_11U_2_else_and_tmp;
  assign m_row2_1_FpMantRNE_23U_11U_2_else_and_tmp = FpMantRNE_23U_11U_2_else_carry_1_sva
      & (FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_2_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1[23]));
  assign m_row1_4_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_sva
      & (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1[23]));
  assign FpMantRNE_23U_11U_1_else_carry_sva = (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_1_mux_73_itm);
  assign FpAdd_6U_10U_1_and_24_ssc = (~(FpAdd_6U_10U_1_and_10_tmp | FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_6_m1c;
  assign FpAdd_6U_10U_1_and_17_ssc = FpAdd_6U_10U_1_and_10_tmp & (~ FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_6_m1c;
  assign FpAdd_6U_10U_1_and_25_ssc = FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_6_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_6_m1c = ~(IsNaN_6U_10U_3_land_3_lpi_1_dfm_3
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_3);
  assign FpAdd_6U_10U_1_and_10_tmp = m_row1_3_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1
      & m_row1_3_FpMantRNE_23U_11U_1_else_and_tmp;
  assign m_row1_3_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_3_sva
      & (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_1_and_22_ssc = (~(FpAdd_6U_10U_1_and_9_tmp | FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_5_m1c;
  assign FpAdd_6U_10U_1_and_15_ssc = FpAdd_6U_10U_1_and_9_tmp & (~ FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_5_m1c;
  assign FpAdd_6U_10U_1_and_23_ssc = FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_5_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_5_m1c = ~(IsNaN_6U_10U_3_land_2_lpi_1_dfm_3
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_3);
  assign FpAdd_6U_10U_1_and_9_tmp = m_row1_2_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1
      & m_row1_2_FpMantRNE_23U_11U_1_else_and_tmp;
  assign m_row1_2_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_2_sva
      & (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_1_and_20_ssc = (~(FpAdd_6U_10U_1_and_8_tmp | FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_4_m1c;
  assign FpAdd_6U_10U_1_and_13_ssc = FpAdd_6U_10U_1_and_8_tmp & (~ FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_4_m1c;
  assign FpAdd_6U_10U_1_and_21_ssc = FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_4_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_4_m1c = ~(IsNaN_6U_10U_3_land_1_lpi_1_dfm_3
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_3);
  assign FpAdd_6U_10U_1_and_8_tmp = m_row1_1_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1
      & m_row1_1_FpMantRNE_23U_11U_1_else_and_tmp;
  assign m_row1_1_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_1_sva
      & (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1[23]));
  assign m_row0_4_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_sva
      & (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1[23]));
  assign FpMantRNE_23U_11U_else_carry_sva = (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1[22:1]), FpAdd_6U_10U_mux_69_itm);
  assign FpAdd_6U_10U_and_24_ssc = (~(FpAdd_6U_10U_and_10_tmp | FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_6_m1c;
  assign FpAdd_6U_10U_and_17_ssc = FpAdd_6U_10U_and_10_tmp & (~ FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_6_m1c;
  assign FpAdd_6U_10U_and_25_ssc = FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_6_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_6_m1c = ~(IsNaN_6U_10U_1_land_3_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_and_10_tmp = m_row0_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 &
      m_row0_3_FpMantRNE_23U_11U_else_and_tmp;
  assign m_row0_3_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_3_sva
      & (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_and_22_ssc = (~(FpAdd_6U_10U_and_9_tmp | FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_and_15_ssc = FpAdd_6U_10U_and_9_tmp & (~ FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_and_23_ssc = FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c = ~(IsNaN_6U_10U_1_land_2_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_and_9_tmp = m_row0_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 & m_row0_2_FpMantRNE_23U_11U_else_and_tmp;
  assign m_row0_2_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_2_sva
      & (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_and_20_ssc = (~(FpAdd_6U_10U_and_8_tmp | FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_4_m1c;
  assign FpAdd_6U_10U_and_13_ssc = FpAdd_6U_10U_and_8_tmp & (~ FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_4_m1c;
  assign FpAdd_6U_10U_and_21_ssc = FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_4_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_4_m1c = ~(IsNaN_6U_10U_1_land_1_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse);
  assign FpAdd_6U_10U_and_8_tmp = m_row0_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 & m_row0_1_FpMantRNE_23U_11U_else_and_tmp;
  assign m_row0_1_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_1_sva
      & (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1[23]));
  assign FpAdd_6U_10U_7_is_a_greater_lor_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_itm_10_1)
      & o_col3_4_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_7_is_a_greater_acc_3_itm_6_1;
  assign nl_FpAdd_6U_10U_7_is_a_greater_acc_3_nl = ({1'b1 , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_7_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_7_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_7_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_7_is_a_greater_acc_3_nl));
  assign FpAdd_6U_10U_7_is_a_greater_lor_3_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_itm_10_1)
      & o_col3_3_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_7_is_a_greater_acc_2_itm_6_1;
  assign nl_FpAdd_6U_10U_7_is_a_greater_acc_2_nl = ({1'b1 , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_7_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_7_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_7_is_a_greater_acc_2_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_7_is_a_greater_acc_2_nl));
  assign FpAdd_6U_10U_7_is_a_greater_lor_2_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_itm_10_1)
      & o_col3_2_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_7_is_a_greater_acc_1_itm_6_1;
  assign nl_FpAdd_6U_10U_7_is_a_greater_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_7_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_7_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_7_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_7_is_a_greater_acc_1_nl));
  assign FpAdd_6U_10U_7_is_a_greater_lor_1_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_itm_10_1)
      & o_col3_1_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_7_is_a_greater_acc_itm_6_1;
  assign nl_FpAdd_6U_10U_7_is_a_greater_acc_nl = ({1'b1 , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_7_is_a_greater_acc_nl = nl_FpAdd_6U_10U_7_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_7_is_a_greater_acc_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_7_is_a_greater_acc_nl));
  assign FpAdd_6U_10U_6_is_a_greater_lor_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_itm_10_1)
      & o_col2_4_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_acc_3_itm_6_1;
  assign nl_FpAdd_6U_10U_6_is_a_greater_acc_3_nl = ({1'b1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_6_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_6_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_6_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_6_is_a_greater_acc_3_nl));
  assign FpAdd_6U_10U_6_is_a_greater_lor_3_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_itm_10_1)
      & o_col2_3_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_acc_2_itm_6_1;
  assign nl_FpAdd_6U_10U_6_is_a_greater_acc_2_nl = ({1'b1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_6_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_6_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_6_is_a_greater_acc_2_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_6_is_a_greater_acc_2_nl));
  assign FpAdd_6U_10U_6_is_a_greater_lor_2_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_itm_10_1)
      & o_col2_2_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_acc_1_itm_6_1;
  assign nl_FpAdd_6U_10U_6_is_a_greater_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_6_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_6_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_6_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_6_is_a_greater_acc_1_nl));
  assign FpAdd_6U_10U_6_is_a_greater_lor_1_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_itm_10_1)
      & o_col2_1_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_acc_itm_6_1;
  assign nl_FpAdd_6U_10U_6_is_a_greater_acc_nl = ({1'b1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_6_is_a_greater_acc_nl = nl_FpAdd_6U_10U_6_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_6_is_a_greater_acc_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_6_is_a_greater_acc_nl));
  assign FpAdd_6U_10U_5_is_a_greater_lor_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_itm_10_1)
      & o_col1_4_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_acc_3_itm_6_1;
  assign nl_FpAdd_6U_10U_5_is_a_greater_acc_3_nl = ({1'b1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_5_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_5_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_5_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_5_is_a_greater_acc_3_nl));
  assign FpAdd_6U_10U_5_is_a_greater_lor_3_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_itm_10_1)
      & o_col1_3_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_acc_2_itm_6_1;
  assign nl_FpAdd_6U_10U_5_is_a_greater_acc_2_nl = ({1'b1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_5_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_5_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_5_is_a_greater_acc_2_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_5_is_a_greater_acc_2_nl));
  assign FpAdd_6U_10U_5_is_a_greater_lor_2_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_itm_10_1)
      & o_col1_2_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_acc_1_itm_6_1;
  assign nl_FpAdd_6U_10U_5_is_a_greater_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_5_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_5_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_5_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_5_is_a_greater_acc_1_nl));
  assign FpAdd_6U_10U_5_is_a_greater_lor_1_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_itm_10_1)
      & o_col1_1_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_acc_itm_6_1;
  assign nl_FpAdd_6U_10U_5_is_a_greater_acc_nl = ({1'b1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_5_is_a_greater_acc_nl = nl_FpAdd_6U_10U_5_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_5_is_a_greater_acc_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_5_is_a_greater_acc_nl));
  assign FpAdd_6U_10U_4_is_a_greater_lor_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_itm_10_1)
      & o_col0_4_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_4_is_a_greater_acc_3_itm_6_1;
  assign nl_FpAdd_6U_10U_4_is_a_greater_acc_3_nl = ({1'b1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_4_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_4_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_4_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_4_is_a_greater_acc_3_nl));
  assign FpAdd_6U_10U_4_is_a_greater_lor_3_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_itm_10_1)
      & o_col0_3_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_4_is_a_greater_acc_2_itm_6_1;
  assign nl_FpAdd_6U_10U_4_is_a_greater_acc_2_nl = ({1'b1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_4_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_4_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_4_is_a_greater_acc_2_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_4_is_a_greater_acc_2_nl));
  assign FpAdd_6U_10U_4_is_a_greater_lor_2_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_itm_10_1)
      & o_col0_2_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_4_is_a_greater_acc_1_itm_6_1;
  assign nl_FpAdd_6U_10U_4_is_a_greater_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_4_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_4_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_4_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_4_is_a_greater_acc_1_nl));
  assign FpAdd_6U_10U_4_is_a_greater_lor_1_lpi_1_dfm_1 = ((~ FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_itm_10_1)
      & o_col0_1_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_4_is_a_greater_acc_itm_6_1;
  assign nl_FpAdd_6U_10U_4_is_a_greater_acc_nl = ({1'b1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2})
      + conv_u2u_6_7({(~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2)}) + 7'b1;
  assign FpAdd_6U_10U_4_is_a_greater_acc_nl = nl_FpAdd_6U_10U_4_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_4_is_a_greater_acc_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_4_is_a_greater_acc_nl));
  assign nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl = nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl[5:0];
  assign o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col0_1_FpNormalize_6U_23U_4_else_lshift_itm, FpNormalize_6U_23U_4_oelse_not_9);
  assign nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl = nl_o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl[5:0];
  assign o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_nl));
  assign nl_o_col0_1_FpNormalize_6U_23U_4_else_acc_nl = ({reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_48)})
      + 6'b1;
  assign o_col0_1_FpNormalize_6U_23U_4_else_acc_nl = nl_o_col0_1_FpNormalize_6U_23U_4_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_nl = MUX_v_6_2_2(6'b000000,
      (o_col0_1_FpNormalize_6U_23U_4_else_acc_nl), FpNormalize_6U_23U_4_oelse_not_9);
  assign nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl = nl_o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_4_nl = (~ o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_4_and_5_nl = o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_nl),
      ({reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2}), (o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23])) , (FpAdd_6U_10U_4_and_4_nl) ,
      (FpAdd_6U_10U_4_and_5_nl)});
  assign nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl = nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl[5:0];
  assign o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col0_2_FpNormalize_6U_23U_4_else_lshift_itm, FpNormalize_6U_23U_4_oelse_not_11);
  assign nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl = nl_o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl[5:0];
  assign o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_nl));
  assign nl_o_col0_2_FpNormalize_6U_23U_4_else_acc_nl = ({reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_49)})
      + 6'b1;
  assign o_col0_2_FpNormalize_6U_23U_4_else_acc_nl = nl_o_col0_2_FpNormalize_6U_23U_4_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_2_nl = MUX_v_6_2_2(6'b000000,
      (o_col0_2_FpNormalize_6U_23U_4_else_acc_nl), FpNormalize_6U_23U_4_oelse_not_11);
  assign nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl = nl_o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_10_nl = (~ o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_4_and_11_nl = o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_2_nl),
      ({reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2}), (o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23])) , (FpAdd_6U_10U_4_and_10_nl)
      , (FpAdd_6U_10U_4_and_11_nl)});
  assign nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl = nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl[5:0];
  assign o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col0_3_FpNormalize_6U_23U_4_else_lshift_itm, FpNormalize_6U_23U_4_oelse_not_13);
  assign nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl = nl_o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl[5:0];
  assign o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_nl));
  assign nl_o_col0_3_FpNormalize_6U_23U_4_else_acc_nl = ({reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_50)})
      + 6'b1;
  assign o_col0_3_FpNormalize_6U_23U_4_else_acc_nl = nl_o_col0_3_FpNormalize_6U_23U_4_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_4_nl = MUX_v_6_2_2(6'b000000,
      (o_col0_3_FpNormalize_6U_23U_4_else_acc_nl), FpNormalize_6U_23U_4_oelse_not_13);
  assign nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl = nl_o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_16_nl = (~ o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_4_and_17_nl = o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_4_nl),
      ({reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2}), (o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23])) , (FpAdd_6U_10U_4_and_16_nl)
      , (FpAdd_6U_10U_4_and_17_nl)});
  assign nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl = nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl[5:0];
  assign o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col0_4_FpNormalize_6U_23U_4_else_lshift_itm, FpNormalize_6U_23U_4_oelse_not_15);
  assign nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_4_o_expo_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl = nl_o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl[5:0];
  assign o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_nl));
  assign nl_o_col0_4_FpNormalize_6U_23U_4_else_acc_nl = ({reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_51)})
      + 6'b1;
  assign o_col0_4_FpNormalize_6U_23U_4_else_acc_nl = nl_o_col0_4_FpNormalize_6U_23U_4_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_6_nl = MUX_v_6_2_2(6'b000000,
      (o_col0_4_FpNormalize_6U_23U_4_else_acc_nl), FpNormalize_6U_23U_4_oelse_not_15);
  assign nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl = nl_o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_4_and_22_nl = (~ o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_4_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_4_and_23_nl = o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_4_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_4_o_expo_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_4_FpNormalize_6U_23U_4_and_6_nl),
      ({reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2}), (o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_4_int_mant_p1_sva_3[23])) , (FpAdd_6U_10U_4_and_22_nl) ,
      (FpAdd_6U_10U_4_and_23_nl)});
  assign nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl = nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl[5:0];
  assign o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col1_1_FpNormalize_6U_23U_5_else_lshift_itm, FpNormalize_6U_23U_5_oelse_not_9);
  assign nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl = nl_o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl[5:0];
  assign o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_nl));
  assign nl_o_col1_1_FpNormalize_6U_23U_5_else_acc_nl = ({reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_52)})
      + 6'b1;
  assign o_col1_1_FpNormalize_6U_23U_5_else_acc_nl = nl_o_col1_1_FpNormalize_6U_23U_5_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_nl = MUX_v_6_2_2(6'b000000,
      (o_col1_1_FpNormalize_6U_23U_5_else_acc_nl), FpNormalize_6U_23U_5_oelse_not_9);
  assign nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl = nl_o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_4_nl = (~ o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_5_and_5_nl = o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_nl),
      ({reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2}), (o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23])) , (FpAdd_6U_10U_5_and_4_nl) ,
      (FpAdd_6U_10U_5_and_5_nl)});
  assign nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl = nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl[5:0];
  assign o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col1_2_FpNormalize_6U_23U_5_else_lshift_itm, FpNormalize_6U_23U_5_oelse_not_11);
  assign nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl = nl_o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl[5:0];
  assign o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_nl));
  assign nl_o_col1_2_FpNormalize_6U_23U_5_else_acc_nl = ({reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_53)})
      + 6'b1;
  assign o_col1_2_FpNormalize_6U_23U_5_else_acc_nl = nl_o_col1_2_FpNormalize_6U_23U_5_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_2_nl = MUX_v_6_2_2(6'b000000,
      (o_col1_2_FpNormalize_6U_23U_5_else_acc_nl), FpNormalize_6U_23U_5_oelse_not_11);
  assign nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl = nl_o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_10_nl = (~ o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_5_and_11_nl = o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_2_nl),
      ({reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2}), (o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23])) , (FpAdd_6U_10U_5_and_10_nl)
      , (FpAdd_6U_10U_5_and_11_nl)});
  assign nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl = nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl[5:0];
  assign o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col1_3_FpNormalize_6U_23U_5_else_lshift_itm, FpNormalize_6U_23U_5_oelse_not_13);
  assign nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl = nl_o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl[5:0];
  assign o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_nl));
  assign nl_o_col1_3_FpNormalize_6U_23U_5_else_acc_nl = ({reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_54)})
      + 6'b1;
  assign o_col1_3_FpNormalize_6U_23U_5_else_acc_nl = nl_o_col1_3_FpNormalize_6U_23U_5_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_4_nl = MUX_v_6_2_2(6'b000000,
      (o_col1_3_FpNormalize_6U_23U_5_else_acc_nl), FpNormalize_6U_23U_5_oelse_not_13);
  assign nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl = nl_o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_16_nl = (~ o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_5_and_17_nl = o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_4_nl),
      ({reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2}), (o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23])) , (FpAdd_6U_10U_5_and_16_nl)
      , (FpAdd_6U_10U_5_and_17_nl)});
  assign nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl = nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl[5:0];
  assign o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col1_4_FpNormalize_6U_23U_5_else_lshift_itm, FpNormalize_6U_23U_5_oelse_not_15);
  assign nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_5_o_expo_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl = nl_o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl[5:0];
  assign o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_nl));
  assign nl_o_col1_4_FpNormalize_6U_23U_5_else_acc_nl = ({reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_55)})
      + 6'b1;
  assign o_col1_4_FpNormalize_6U_23U_5_else_acc_nl = nl_o_col1_4_FpNormalize_6U_23U_5_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_6_nl = MUX_v_6_2_2(6'b000000,
      (o_col1_4_FpNormalize_6U_23U_5_else_acc_nl), FpNormalize_6U_23U_5_oelse_not_15);
  assign nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl = nl_o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_5_and_22_nl = (~ o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_5_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_5_and_23_nl = o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_5_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_5_o_expo_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_5_FpNormalize_6U_23U_5_and_6_nl),
      ({reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2}), (o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_5_int_mant_p1_sva_3[23])) , (FpAdd_6U_10U_5_and_22_nl) ,
      (FpAdd_6U_10U_5_and_23_nl)});
  assign nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl = nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl[5:0];
  assign o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col2_1_FpNormalize_6U_23U_6_else_lshift_itm, FpNormalize_6U_23U_6_oelse_not_9);
  assign nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl = nl_o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl[5:0];
  assign o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_nl));
  assign nl_o_col2_1_FpNormalize_6U_23U_6_else_acc_nl = ({reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_56)})
      + 6'b1;
  assign o_col2_1_FpNormalize_6U_23U_6_else_acc_nl = nl_o_col2_1_FpNormalize_6U_23U_6_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_nl = MUX_v_6_2_2(6'b000000,
      (o_col2_1_FpNormalize_6U_23U_6_else_acc_nl), FpNormalize_6U_23U_6_oelse_not_9);
  assign nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl = nl_o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_4_nl = (~ o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_6_and_5_nl = o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_nl),
      ({reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2}), (o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23])) , (FpAdd_6U_10U_6_and_4_nl) ,
      (FpAdd_6U_10U_6_and_5_nl)});
  assign nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl = nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl[5:0];
  assign o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col2_2_FpNormalize_6U_23U_6_else_lshift_itm, FpNormalize_6U_23U_6_oelse_not_11);
  assign nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl = nl_o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl[5:0];
  assign o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_nl));
  assign nl_o_col2_2_FpNormalize_6U_23U_6_else_acc_nl = ({reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_57)})
      + 6'b1;
  assign o_col2_2_FpNormalize_6U_23U_6_else_acc_nl = nl_o_col2_2_FpNormalize_6U_23U_6_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_2_nl = MUX_v_6_2_2(6'b000000,
      (o_col2_2_FpNormalize_6U_23U_6_else_acc_nl), FpNormalize_6U_23U_6_oelse_not_11);
  assign nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl = nl_o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_10_nl = (~ o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_6_and_11_nl = o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_2_nl),
      ({reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2}), (o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23])) , (FpAdd_6U_10U_6_and_10_nl)
      , (FpAdd_6U_10U_6_and_11_nl)});
  assign nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl = nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl[5:0];
  assign o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col2_3_FpNormalize_6U_23U_6_else_lshift_itm, FpNormalize_6U_23U_6_oelse_not_13);
  assign nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl = nl_o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl[5:0];
  assign o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_nl));
  assign nl_o_col2_3_FpNormalize_6U_23U_6_else_acc_nl = ({reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_58)})
      + 6'b1;
  assign o_col2_3_FpNormalize_6U_23U_6_else_acc_nl = nl_o_col2_3_FpNormalize_6U_23U_6_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_4_nl = MUX_v_6_2_2(6'b000000,
      (o_col2_3_FpNormalize_6U_23U_6_else_acc_nl), FpNormalize_6U_23U_6_oelse_not_13);
  assign nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl = nl_o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_16_nl = (~ o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_6_and_17_nl = o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_4_nl),
      ({reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2}), (o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23])) , (FpAdd_6U_10U_6_and_16_nl)
      , (FpAdd_6U_10U_6_and_17_nl)});
  assign nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl = nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl[5:0];
  assign o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col2_4_FpNormalize_6U_23U_6_else_lshift_itm, FpNormalize_6U_23U_6_oelse_not_15);
  assign nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_6_o_expo_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl = nl_o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl[5:0];
  assign o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_nl));
  assign nl_o_col2_4_FpNormalize_6U_23U_6_else_acc_nl = ({reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_59)})
      + 6'b1;
  assign o_col2_4_FpNormalize_6U_23U_6_else_acc_nl = nl_o_col2_4_FpNormalize_6U_23U_6_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_6_nl = MUX_v_6_2_2(6'b000000,
      (o_col2_4_FpNormalize_6U_23U_6_else_acc_nl), FpNormalize_6U_23U_6_oelse_not_15);
  assign nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl = nl_o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_6_and_22_nl = (~ o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_6_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_6_and_23_nl = o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_6_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_6_o_expo_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_6_FpNormalize_6U_23U_6_and_6_nl),
      ({reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2}), (o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_6_int_mant_p1_sva_3[23])) , (FpAdd_6U_10U_6_and_22_nl) ,
      (FpAdd_6U_10U_6_and_23_nl)});
  assign nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl = nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl[5:0];
  assign o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col3_1_FpNormalize_6U_23U_7_else_lshift_itm, FpNormalize_6U_23U_7_oelse_not_9);
  assign nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl = nl_o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl[5:0];
  assign o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_nl));
  assign nl_o_col3_1_FpNormalize_6U_23U_7_else_acc_nl = ({reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_60)})
      + 6'b1;
  assign o_col3_1_FpNormalize_6U_23U_7_else_acc_nl = nl_o_col3_1_FpNormalize_6U_23U_7_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_nl = MUX_v_6_2_2(6'b000000,
      (o_col3_1_FpNormalize_6U_23U_7_else_acc_nl), FpNormalize_6U_23U_7_oelse_not_9);
  assign nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl = nl_o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_4_nl = (~ o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_7_and_5_nl = o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23]);
  assign FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_nl),
      ({reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2}), (o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23])) , (FpAdd_6U_10U_7_and_4_nl) ,
      (FpAdd_6U_10U_7_and_5_nl)});
  assign nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl = nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl[5:0];
  assign o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col3_2_FpNormalize_6U_23U_7_else_lshift_itm, FpNormalize_6U_23U_7_oelse_not_11);
  assign nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl = nl_o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl[5:0];
  assign o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_nl));
  assign nl_o_col3_2_FpNormalize_6U_23U_7_else_acc_nl = ({reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_61)})
      + 6'b1;
  assign o_col3_2_FpNormalize_6U_23U_7_else_acc_nl = nl_o_col3_2_FpNormalize_6U_23U_7_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_2_nl = MUX_v_6_2_2(6'b000000,
      (o_col3_2_FpNormalize_6U_23U_7_else_acc_nl), FpNormalize_6U_23U_7_oelse_not_11);
  assign nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl = nl_o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_10_nl = (~ o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_7_and_11_nl = o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23]);
  assign FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_2_nl),
      ({reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2}), (o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23])) , (FpAdd_6U_10U_7_and_10_nl)
      , (FpAdd_6U_10U_7_and_11_nl)});
  assign nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl = nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl[5:0];
  assign o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col3_3_FpNormalize_6U_23U_7_else_lshift_itm, FpNormalize_6U_23U_7_oelse_not_13);
  assign nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl = nl_o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl[5:0];
  assign o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_nl));
  assign nl_o_col3_3_FpNormalize_6U_23U_7_else_acc_nl = ({reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_62)})
      + 6'b1;
  assign o_col3_3_FpNormalize_6U_23U_7_else_acc_nl = nl_o_col3_3_FpNormalize_6U_23U_7_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_4_nl = MUX_v_6_2_2(6'b000000,
      (o_col3_3_FpNormalize_6U_23U_7_else_acc_nl), FpNormalize_6U_23U_7_oelse_not_13);
  assign nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl = nl_o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_16_nl = (~ o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_7_and_17_nl = o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23]);
  assign FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_4_nl),
      ({reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2}), (o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23])) , (FpAdd_6U_10U_7_and_16_nl)
      , (FpAdd_6U_10U_7_and_17_nl)});
  assign nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1 , (reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2[3:1])})
      + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl = nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl[5:0];
  assign o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      o_col3_4_FpNormalize_6U_23U_7_else_lshift_itm, FpNormalize_6U_23U_7_oelse_not_15);
  assign nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_7_o_expo_lpi_1_dfm_2[5:1])})
      + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl = nl_o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl[5:0];
  assign o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_nl));
  assign nl_o_col3_4_FpNormalize_6U_23U_7_else_acc_nl = ({reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2})
      + ({1'b1 , (~ libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_63)})
      + 6'b1;
  assign o_col3_4_FpNormalize_6U_23U_7_else_acc_nl = nl_o_col3_4_FpNormalize_6U_23U_7_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_6_nl = MUX_v_6_2_2(6'b000000,
      (o_col3_4_FpNormalize_6U_23U_7_else_acc_nl), FpNormalize_6U_23U_7_oelse_not_15);
  assign nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl = ({reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp
      , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1 , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2})
      + 6'b1;
  assign o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl = nl_o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl[5:0];
  assign FpAdd_6U_10U_7_and_22_nl = (~ o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_7_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_7_and_23_nl = o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_7_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_7_o_expo_lpi_1_dfm_2 = MUX1HOT_v_6_3_2((FpNormalize_6U_23U_7_FpNormalize_6U_23U_7_and_6_nl),
      ({reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1
      , reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2}), (o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_nl),
      {(~ (FpAdd_6U_10U_7_int_mant_p1_sva_3[23])) , (FpAdd_6U_10U_7_and_22_nl) ,
      (FpAdd_6U_10U_7_and_23_nl)});
  assign o_col3_4_FpMantRNE_23U_11U_7_else_and_tmp = FpMantRNE_23U_11U_7_else_carry_sva
      & (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_7_int_mant_p1_sva_3[23]));
  assign FpMantRNE_23U_11U_7_else_carry_sva = (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_7_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_7_int_mant_p1_sva_3[22:1]), FpAdd_6U_10U_7_int_mant_p1_sva_3[23]);
  assign o_col3_3_FpMantRNE_23U_11U_7_else_and_tmp = FpMantRNE_23U_11U_7_else_carry_3_sva
      & (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23]));
  assign FpMantRNE_23U_11U_7_else_carry_3_sva = (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_7_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[22:1]), FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23]);
  assign o_col3_2_FpMantRNE_23U_11U_7_else_and_tmp = FpMantRNE_23U_11U_7_else_carry_2_sva
      & (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23]));
  assign FpMantRNE_23U_11U_7_else_carry_2_sva = (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_7_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[22:1]), FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23]);
  assign o_col3_1_FpMantRNE_23U_11U_7_else_and_tmp = FpMantRNE_23U_11U_7_else_carry_1_sva
      & (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23]));
  assign FpMantRNE_23U_11U_7_else_carry_1_sva = (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_7_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[22:1]), FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23]);
  assign o_col2_4_FpMantRNE_23U_11U_6_else_and_tmp = FpMantRNE_23U_11U_6_else_carry_sva
      & (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_6_int_mant_p1_sva_3[23]));
  assign FpMantRNE_23U_11U_6_else_carry_sva = (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_6_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_6_int_mant_p1_sva_3[22:1]), FpAdd_6U_10U_6_int_mant_p1_sva_3[23]);
  assign o_col2_3_FpMantRNE_23U_11U_6_else_and_tmp = FpMantRNE_23U_11U_6_else_carry_3_sva
      & (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23]));
  assign FpMantRNE_23U_11U_6_else_carry_3_sva = (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_6_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[22:1]), FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23]);
  assign o_col2_2_FpMantRNE_23U_11U_6_else_and_tmp = FpMantRNE_23U_11U_6_else_carry_2_sva
      & (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23]));
  assign FpMantRNE_23U_11U_6_else_carry_2_sva = (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_6_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[22:1]), FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23]);
  assign o_col2_1_FpMantRNE_23U_11U_6_else_and_tmp = FpMantRNE_23U_11U_6_else_carry_1_sva
      & (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23]));
  assign FpMantRNE_23U_11U_6_else_carry_1_sva = (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_6_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[22:1]), FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23]);
  assign o_col1_4_FpMantRNE_23U_11U_5_else_and_tmp = FpMantRNE_23U_11U_5_else_carry_sva
      & (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_5_int_mant_p1_sva_3[23]));
  assign FpMantRNE_23U_11U_5_else_carry_sva = (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_5_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_5_int_mant_p1_sva_3[22:1]), FpAdd_6U_10U_5_int_mant_p1_sva_3[23]);
  assign o_col1_3_FpMantRNE_23U_11U_5_else_and_tmp = FpMantRNE_23U_11U_5_else_carry_3_sva
      & (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23]));
  assign FpMantRNE_23U_11U_5_else_carry_3_sva = (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_5_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[22:1]), FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23]);
  assign o_col1_2_FpMantRNE_23U_11U_5_else_and_tmp = FpMantRNE_23U_11U_5_else_carry_2_sva
      & (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23]));
  assign FpMantRNE_23U_11U_5_else_carry_2_sva = (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_5_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[22:1]), FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23]);
  assign o_col1_1_FpMantRNE_23U_11U_5_else_and_tmp = FpMantRNE_23U_11U_5_else_carry_1_sva
      & (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23]));
  assign FpMantRNE_23U_11U_5_else_carry_1_sva = (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_5_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[22:1]), FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23]);
  assign o_col0_4_FpMantRNE_23U_11U_4_else_and_tmp = FpMantRNE_23U_11U_4_else_carry_sva
      & (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_4_int_mant_p1_sva_3[23]));
  assign FpMantRNE_23U_11U_4_else_carry_sva = (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_4_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_4_int_mant_p1_sva_3[22:1]), FpAdd_6U_10U_4_int_mant_p1_sva_3[23]);
  assign o_col0_3_FpMantRNE_23U_11U_4_else_and_tmp = FpMantRNE_23U_11U_4_else_carry_3_sva
      & (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23]));
  assign FpMantRNE_23U_11U_4_else_carry_3_sva = (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_4_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[22:1]), FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23]);
  assign o_col0_2_FpMantRNE_23U_11U_4_else_and_tmp = FpMantRNE_23U_11U_4_else_carry_2_sva
      & (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23]));
  assign FpMantRNE_23U_11U_4_else_carry_2_sva = (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_4_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[22:1]), FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23]);
  assign o_col0_1_FpMantRNE_23U_11U_4_else_and_tmp = FpMantRNE_23U_11U_4_else_carry_1_sva
      & (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23]));
  assign FpMantRNE_23U_11U_4_else_carry_1_sva = (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_4_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[22:1]), FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23]);
  assign IsNaN_6U_10U_16_land_lpi_1_dfm = ~(IsNaN_6U_10U_16_nor_15_itm_2 | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_165_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva[9:0]),
      FpAdd_6U_10U_7_o_mant_lpi_2, data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_253_nl = ~ data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_165_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_253_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl),
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_7_o_mant_lpi_2,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_nl),
      or_tmp_510);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_154_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva[9:0]),
      FpAdd_6U_10U_6_o_mant_lpi_2, data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_251_nl = ~ data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_154_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_251_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl),
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_1_nl),
      FpAdd_6U_10U_6_o_mant_lpi_2, IsNaN_6U_10U_16_land_15_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_143_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva[9:0]),
      FpAdd_6U_10U_5_o_mant_lpi_2, data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_249_nl = ~ data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_143_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_249_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl),
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_2_nl),
      FpAdd_6U_10U_5_o_mant_lpi_2, IsNaN_6U_10U_16_land_14_lpi_1_dfm_3);
  assign IsNaN_6U_10U_16_land_13_lpi_1_dfm = ~(IsNaN_6U_10U_16_nor_12_itm_2 | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_132_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva[9:0]),
      FpAdd_6U_10U_4_o_mant_lpi_2, data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_247_nl = ~ data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_132_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_247_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl),
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_3_mx0 = MUX_v_10_2_2(FpAdd_6U_10U_4_o_mant_lpi_2,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_3_nl),
      or_tmp_576);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_121_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva[9:0]),
      FpAdd_6U_10U_7_o_mant_3_lpi_2, data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_245_nl = ~ data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_121_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_245_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl),
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_4_nl),
      FpAdd_6U_10U_7_o_mant_3_lpi_2, IsNaN_6U_10U_16_land_12_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_110_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva[9:0]),
      FpAdd_6U_10U_6_o_mant_3_lpi_2, data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_243_nl = ~ data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_110_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_243_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl),
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_5_nl),
      FpAdd_6U_10U_6_o_mant_3_lpi_2, IsNaN_6U_10U_16_land_11_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_99_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva[9:0]),
      FpAdd_6U_10U_5_o_mant_3_lpi_2, data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_241_nl = ~ data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_99_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_241_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl),
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_6_nl),
      FpAdd_6U_10U_5_o_mant_3_lpi_2, IsNaN_6U_10U_16_land_10_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_88_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva[9:0]),
      FpAdd_6U_10U_4_o_mant_3_lpi_2, data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_239_nl = ~ data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_88_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_239_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl),
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_7_nl),
      FpAdd_6U_10U_4_o_mant_3_lpi_2, IsNaN_6U_10U_16_land_9_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_77_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva[9:0]),
      FpAdd_6U_10U_7_o_mant_2_lpi_2, data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_237_nl = ~ data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_77_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_237_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl),
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_8_nl),
      FpAdd_6U_10U_7_o_mant_2_lpi_2, IsNaN_6U_10U_16_land_8_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_66_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva[9:0]),
      FpAdd_6U_10U_6_o_mant_2_lpi_2, data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_235_nl = ~ data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_66_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_235_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl),
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_9_nl),
      FpAdd_6U_10U_6_o_mant_2_lpi_2, IsNaN_6U_10U_16_land_7_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_55_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva[9:0]),
      FpAdd_6U_10U_5_o_mant_2_lpi_2, data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_233_nl = ~ data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_55_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_233_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl),
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_10_nl),
      FpAdd_6U_10U_5_o_mant_2_lpi_2, IsNaN_6U_10U_16_land_6_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_44_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva[9:0]),
      FpAdd_6U_10U_4_o_mant_2_lpi_2, data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_231_nl = ~ data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_44_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_231_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl),
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_11_nl),
      FpAdd_6U_10U_4_o_mant_2_lpi_2, IsNaN_6U_10U_16_land_5_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_33_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva[9:0]),
      FpAdd_6U_10U_7_o_mant_1_lpi_2, data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_229_nl = ~ data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_33_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_229_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl),
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_12_nl),
      FpAdd_6U_10U_7_o_mant_1_lpi_2, IsNaN_6U_10U_16_land_4_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_22_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva[9:0]),
      FpAdd_6U_10U_6_o_mant_1_lpi_2, data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_227_nl = ~ data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_22_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_227_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl),
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_13_nl),
      FpAdd_6U_10U_6_o_mant_1_lpi_2, IsNaN_6U_10U_16_land_3_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_11_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva[9:0]),
      FpAdd_6U_10U_5_o_mant_1_lpi_2, data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_225_nl = ~ data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_11_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_225_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl),
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_14_nl),
      FpAdd_6U_10U_5_o_mant_1_lpi_2, IsNaN_6U_10U_16_land_2_lpi_1_dfm_3);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_nl = MUX_v_10_2_2((FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva[9:0]),
      FpAdd_6U_10U_4_o_mant_1_lpi_2, data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_223_nl = ~ data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl = ~(MUX_v_10_2_2(10'b0000000000,
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_nl), (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_223_nl)));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl
      = ~(MUX_v_10_2_2(10'b0000000000, (FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl),
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_FpExpoWidthDec_6U_5U_10U_1U_1U_nand_15_nl),
      FpAdd_6U_10U_4_o_mant_1_lpi_2, IsNaN_6U_10U_16_land_1_lpi_1_dfm_3);
  assign data_truncate_1_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_1_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_1_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_1_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_1_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_1_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva = data_truncate_1_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_1_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva
      = (~ (FpAdd_6U_10U_4_o_expo_1_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_2_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_1_sva = FpAdd_6U_10U_4_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_1_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_1_sva = FpAdd_6U_10U_4_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_1_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_1_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_1_sva = FpAdd_6U_10U_4_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_1_sva[9:0]);
  assign data_truncate_2_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_2_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_2_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_2_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_2_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_2_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva = data_truncate_2_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_2_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva
      = (~ (FpAdd_6U_10U_5_o_expo_1_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_3_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_2_sva = FpAdd_6U_10U_5_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_2_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_2_sva = FpAdd_6U_10U_5_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_2_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_2_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_2_sva = FpAdd_6U_10U_5_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_2_sva[9:0]);
  assign data_truncate_3_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_3_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_3_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_3_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_3_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_3_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva = data_truncate_3_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_3_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva
      = (~ (FpAdd_6U_10U_6_o_expo_1_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_4_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_3_sva = FpAdd_6U_10U_6_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_3_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_3_sva = FpAdd_6U_10U_6_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_3_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_3_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_3_sva = FpAdd_6U_10U_6_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_3_sva[9:0]);
  assign data_truncate_4_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_4_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_4_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_4_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_4_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_4_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva = data_truncate_4_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_4_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva
      = (~ (FpAdd_6U_10U_7_o_expo_1_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_5_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_4_sva = FpAdd_6U_10U_7_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_4_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_4_sva = FpAdd_6U_10U_7_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_4_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_4_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_4_sva = FpAdd_6U_10U_7_o_mant_1_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_4_sva[9:0]);
  assign data_truncate_5_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_5_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_5_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_5_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_5_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_5_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva = data_truncate_5_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_5_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva
      = (~ (FpAdd_6U_10U_4_o_expo_2_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_6_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_5_sva = FpAdd_6U_10U_4_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_5_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_5_sva = FpAdd_6U_10U_4_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_5_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_5_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_5_sva = FpAdd_6U_10U_4_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_5_sva[9:0]);
  assign data_truncate_6_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_6_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_6_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_6_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_6_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_6_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva = data_truncate_6_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_6_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva
      = (~ (FpAdd_6U_10U_5_o_expo_2_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_7_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_6_sva = FpAdd_6U_10U_5_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_6_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_6_sva = FpAdd_6U_10U_5_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_6_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_6_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_6_sva = FpAdd_6U_10U_5_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_6_sva[9:0]);
  assign data_truncate_7_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_7_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_7_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_7_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_7_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_7_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva = data_truncate_7_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_7_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva
      = (~ (FpAdd_6U_10U_6_o_expo_2_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_8_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_7_sva = FpAdd_6U_10U_6_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_7_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_7_sva = FpAdd_6U_10U_6_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_7_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_7_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_7_sva = FpAdd_6U_10U_6_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_7_sva[9:0]);
  assign data_truncate_8_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_8_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_8_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_8_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_8_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_8_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva = data_truncate_8_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_8_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva
      = (~ (FpAdd_6U_10U_7_o_expo_2_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_9_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_8_sva = FpAdd_6U_10U_7_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_8_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_8_sva = FpAdd_6U_10U_7_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_8_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_8_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_8_sva = FpAdd_6U_10U_7_o_mant_2_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_8_sva[9:0]);
  assign data_truncate_9_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_9_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_9_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_9_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_9_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_9_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva = data_truncate_9_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_9_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva
      = (~ (FpAdd_6U_10U_4_o_expo_3_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_10_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_9_sva = FpAdd_6U_10U_4_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_9_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_9_sva = FpAdd_6U_10U_4_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_9_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_9_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_9_sva = FpAdd_6U_10U_4_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_9_sva[9:0]);
  assign data_truncate_10_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_10_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_10_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_10_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_10_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_10_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva = data_truncate_10_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_10_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva
      = (~ (FpAdd_6U_10U_5_o_expo_3_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_11_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_10_sva = FpAdd_6U_10U_5_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_10_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_10_sva = FpAdd_6U_10U_5_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_10_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_10_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_10_sva = FpAdd_6U_10U_5_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_10_sva[9:0]);
  assign data_truncate_11_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_11_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_11_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_11_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_11_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_11_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva = data_truncate_11_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_11_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva
      = (~ (FpAdd_6U_10U_6_o_expo_3_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_12_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_11_sva = FpAdd_6U_10U_6_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_11_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_11_sva = FpAdd_6U_10U_6_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_11_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_11_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_11_sva = FpAdd_6U_10U_6_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_11_sva[9:0]);
  assign data_truncate_12_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_12_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_12_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_12_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_12_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_12_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva = data_truncate_12_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_12_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva
      = (~ (FpAdd_6U_10U_7_o_expo_3_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_13_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_12_sva = FpAdd_6U_10U_7_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_12_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_12_sva = FpAdd_6U_10U_7_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_12_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_12_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_12_sva = FpAdd_6U_10U_7_o_mant_3_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_12_sva[9:0]);
  assign data_truncate_13_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_13_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_13_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_13_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_13_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_13_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva = data_truncate_13_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_13_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva
      = (~ (FpAdd_6U_10U_4_o_expo_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_14_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_13_sva = FpAdd_6U_10U_4_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_13_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_13_sva = FpAdd_6U_10U_4_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_13_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_13_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_13_sva = FpAdd_6U_10U_4_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_13_sva[9:0]);
  assign data_truncate_14_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_14_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_14_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_14_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_14_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_14_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva = data_truncate_14_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_14_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva
      = (~ (FpAdd_6U_10U_5_o_expo_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_15_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_14_sva = FpAdd_6U_10U_5_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_14_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_14_sva = FpAdd_6U_10U_5_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_14_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_14_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_14_sva = FpAdd_6U_10U_5_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_14_sva[9:0]);
  assign data_truncate_15_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_15_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_15_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_15_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_15_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_15_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva = data_truncate_15_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_15_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva
      = (~ (FpAdd_6U_10U_6_o_expo_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva =
      nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_16_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_15_sva = FpAdd_6U_10U_6_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_15_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_15_sva = FpAdd_6U_10U_6_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_15_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_15_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_15_sva = FpAdd_6U_10U_6_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_15_sva[9:0]);
  assign data_truncate_16_FpMantDecShiftRight_10U_6U_10U_carry_and_nl = ((FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_guard_mask_sva[10])) & ((FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_stick_mask_sva[10]) | (FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_sva!=10'b0000000000)
      | (FpMantDecShiftRight_10U_6U_10U_least_mask_sva[10]));
  assign nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva = data_truncate_16_FpMantDecShiftRight_10U_6U_10U_i_mant_s_rshift_itm
      + conv_u2u_1_11(data_truncate_16_FpMantDecShiftRight_10U_6U_10U_carry_and_nl);
  assign FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva = nl_FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva[10:0];
  assign nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva
      = (~ (FpAdd_6U_10U_7_o_expo_lpi_2[3:1])) + 3'b1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva = nl_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_if_i_shift_acc_psp_1_sva[2:0];
  assign FpMantDecShiftRight_10U_6U_10U_guard_bits_9_0_sva = FpAdd_6U_10U_7_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_guard_mask_sva[9:0]);
  assign FpMantDecShiftRight_10U_6U_10U_stick_bits_9_0_sva = FpAdd_6U_10U_7_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_stick_mask_sva[9:0]);
  assign nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_sva = FpMantDecShiftRight_10U_6U_10U_guard_mask_sva
      + 11'b11111111111;
  assign FpMantDecShiftRight_10U_6U_10U_stick_mask_sva = nl_FpMantDecShiftRight_10U_6U_10U_stick_mask_sva[10:0];
  assign FpMantDecShiftRight_10U_6U_10U_least_bits_9_0_sva = FpAdd_6U_10U_7_o_mant_lpi_2
      & (FpMantDecShiftRight_10U_6U_10U_least_mask_sva[9:0]);
  assign main_stage_en_1 = chn_data_in_rsci_bawt & or_181_cse;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_15_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_3_o_expo_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse , FpAdd_6U_10U_3_and_26_ssc
      , FpAdd_6U_10U_3_and_19_ssc});
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_5 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_15_nl)
      | FpAdd_6U_10U_3_and_27_ssc;
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_7,
      FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_3_o_expo_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse , FpAdd_6U_10U_3_and_26_ssc
      , FpAdd_6U_10U_3_and_19_ssc , FpAdd_6U_10U_3_and_27_ssc});
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_3_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_3_o_expo_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse , FpAdd_6U_10U_3_and_26_ssc
      , FpAdd_6U_10U_3_and_19_ssc});
  assign FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_4 = (FpAdd_6U_10U_3_FpAdd_6U_10U_3_mux1h_3_nl)
      | FpAdd_6U_10U_3_and_27_ssc;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_15_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_2_o_expo_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse , FpAdd_6U_10U_2_and_26_ssc
      , FpAdd_6U_10U_2_and_19_ssc});
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_5 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_15_nl)
      | FpAdd_6U_10U_2_and_27_ssc;
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_7,
      FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_2_o_expo_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse , FpAdd_6U_10U_2_and_26_ssc
      , FpAdd_6U_10U_2_and_19_ssc , FpAdd_6U_10U_2_and_27_ssc});
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_3_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_2_o_expo_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse , FpAdd_6U_10U_2_and_26_ssc
      , FpAdd_6U_10U_2_and_19_ssc});
  assign FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_4 = (FpAdd_6U_10U_2_FpAdd_6U_10U_2_mux1h_3_nl)
      | FpAdd_6U_10U_2_and_27_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_15_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_1_o_expo_sva_4[5]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse , FpAdd_6U_10U_1_and_26_ssc
      , FpAdd_6U_10U_1_and_19_ssc});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_15_nl)
      | FpAdd_6U_10U_1_and_27_ssc;
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_7,
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_1_o_expo_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse , FpAdd_6U_10U_1_and_26_ssc
      , FpAdd_6U_10U_1_and_19_ssc , FpAdd_6U_10U_1_and_27_ssc});
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_3_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_1_o_expo_sva_4[4]),
      {FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse , FpAdd_6U_10U_1_and_26_ssc
      , FpAdd_6U_10U_1_and_19_ssc});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_3_nl)
      | FpAdd_6U_10U_1_and_27_ssc;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_1_1,
      FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_mx0, (FpAdd_6U_10U_o_expo_sva_4[5]), {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse
      , FpAdd_6U_10U_and_26_ssc , FpAdd_6U_10U_and_19_ssc});
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl)
      | FpAdd_6U_10U_and_27_ssc;
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_7,
      FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0_mx0, (FpAdd_6U_10U_o_expo_sva_4[3:0]),
      4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse , FpAdd_6U_10U_and_26_ssc
      , FpAdd_6U_10U_and_19_ssc , FpAdd_6U_10U_and_27_ssc});
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_3_nl = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_0_1,
      FpAdd_6U_10U_o_expo_lpi_1_dfm_2_4_mx0, (FpAdd_6U_10U_o_expo_sva_4[4]), {FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse
      , FpAdd_6U_10U_and_26_ssc , FpAdd_6U_10U_and_19_ssc});
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_7_4 = (FpAdd_6U_10U_FpAdd_6U_10U_mux1h_3_nl)
      | FpAdd_6U_10U_and_27_ssc;
  assign nl_FpAdd_6U_10U_o_expo_sva_4 = ({FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_mx0 ,
      FpAdd_6U_10U_o_expo_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_sva_4 = nl_FpAdd_6U_10U_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl = FpAdd_6U_10U_is_inf_lpi_1_dfm
      | (~ m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl), m_row0_4_FpMantRNE_23U_11U_else_and_tmp);
  assign FpAdd_6U_10U_is_inf_lpi_1_dfm = ~(m_row0_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1[23])));
  assign nl_m_row0_4_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_sva);
  assign m_row0_4_FpMantRNE_23U_11U_else_acc_nl = nl_m_row0_4_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_11_itm = MUX_v_10_2_2((m_row0_4_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_1_o_expo_sva_4 = ({FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_sva_4 = nl_FpAdd_6U_10U_1_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl = FpAdd_6U_10U_1_is_inf_lpi_1_dfm
      | (~ m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl), m_row1_4_FpMantRNE_23U_11U_1_else_and_tmp);
  assign FpAdd_6U_10U_1_is_inf_lpi_1_dfm = ~(m_row1_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1[23])));
  assign nl_m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_sva);
  assign m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl = nl_m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_11_itm = MUX_v_10_2_2((m_row1_4_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_2_o_expo_sva_4 = ({FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_2_o_expo_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_2_o_expo_sva_4 = nl_FpAdd_6U_10U_2_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_3_nl = FpAdd_6U_10U_2_is_inf_lpi_1_dfm
      | (~ m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_2_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_2_if_4_FpAdd_6U_10U_2_if_4_or_3_nl), m_row2_4_FpMantRNE_23U_11U_2_else_and_tmp);
  assign FpAdd_6U_10U_2_is_inf_lpi_1_dfm = ~(m_row2_4_FpAdd_6U_10U_2_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1[23])));
  assign nl_m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl = (FpAdd_6U_10U_2_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_2_else_carry_sva);
  assign m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl = nl_m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl[9:0];
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_11_itm = MUX_v_10_2_2((m_row2_4_FpMantRNE_23U_11U_2_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0);
  assign nl_FpAdd_6U_10U_3_o_expo_sva_4 = ({FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_5_mx0
      , FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_4_mx0 , FpAdd_6U_10U_3_o_expo_lpi_1_dfm_2_3_0_mx0})
      + 6'b1;
  assign FpAdd_6U_10U_3_o_expo_sva_4 = nl_FpAdd_6U_10U_3_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_3_nl = FpAdd_6U_10U_3_is_inf_lpi_1_dfm
      | (~ m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_3_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_3_if_4_FpAdd_6U_10U_3_if_4_or_3_nl), m_row3_4_FpMantRNE_23U_11U_3_else_and_tmp);
  assign FpAdd_6U_10U_3_is_inf_lpi_1_dfm = ~(m_row3_4_FpAdd_6U_10U_3_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1[23])));
  assign nl_m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl = (FpAdd_6U_10U_3_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_3_else_carry_sva);
  assign m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl = nl_m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl[9:0];
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_11_itm = MUX_v_10_2_2((m_row3_4_FpMantRNE_23U_11U_3_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0);
  assign FpAdd_6U_10U_3_and_26_ssc = (~(FpAdd_6U_10U_3_and_11_tmp | FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_7_m1c;
  assign FpAdd_6U_10U_3_and_19_ssc = FpAdd_6U_10U_3_and_11_tmp & (~ FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_7_m1c;
  assign FpAdd_6U_10U_3_and_27_ssc = FpAdd_6U_10U_3_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_7_m1c;
  assign FpAdd_6U_10U_3_FpAdd_6U_10U_3_nor_7_m1c = ~(IsNaN_6U_10U_7_land_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse);
  assign FpAdd_6U_10U_3_and_11_tmp = m_row3_4_FpAdd_6U_10U_3_if_4_if_acc_1_itm_5_1
      & m_row3_4_FpMantRNE_23U_11U_3_else_and_tmp;
  assign FpAdd_6U_10U_2_and_26_ssc = (~(FpAdd_6U_10U_2_and_11_tmp | FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_7_m1c;
  assign FpAdd_6U_10U_2_and_19_ssc = FpAdd_6U_10U_2_and_11_tmp & (~ FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_7_m1c;
  assign FpAdd_6U_10U_2_and_27_ssc = FpAdd_6U_10U_2_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_7_m1c;
  assign FpAdd_6U_10U_2_FpAdd_6U_10U_2_nor_7_m1c = ~(IsNaN_6U_10U_5_land_lpi_1_dfm_3
      | IsNaN_6U_10U_4_land_lpi_1_dfm_st_2);
  assign FpAdd_6U_10U_2_and_11_tmp = m_row2_4_FpAdd_6U_10U_2_if_4_if_acc_1_itm_5_1
      & m_row2_4_FpMantRNE_23U_11U_2_else_and_tmp;
  assign FpAdd_6U_10U_1_and_26_ssc = (~(FpAdd_6U_10U_1_and_11_tmp | FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_and_19_ssc = FpAdd_6U_10U_1_and_11_tmp & (~ FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_and_27_ssc = FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c = ~(IsNaN_6U_10U_3_land_lpi_1_dfm_3
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_2);
  assign FpAdd_6U_10U_1_and_11_tmp = m_row1_4_FpAdd_6U_10U_1_if_4_if_acc_1_itm_5_1
      & m_row1_4_FpMantRNE_23U_11U_1_else_and_tmp;
  assign FpAdd_6U_10U_and_26_ssc = (~(FpAdd_6U_10U_and_11_tmp | FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_and_19_ssc = FpAdd_6U_10U_and_11_tmp & (~ FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_and_27_ssc = FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c = ~(IsNaN_6U_10U_1_land_lpi_1_dfm_3
      | reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse);
  assign FpAdd_6U_10U_and_11_tmp = m_row0_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 &
      m_row0_4_FpMantRNE_23U_11U_else_and_tmp;
  assign FpAdd_6U_10U_4_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_a_int_mant_p1_1_sva,
      FpAdd_6U_10U_4_addend_larger_asn_19_mx0w1, and_dcpl_449);
  assign FpAdd_6U_10U_4_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_asn_19_mx0w1,
      FpAdd_6U_10U_4_a_int_mant_p1_1_sva, and_dcpl_449);
  assign FpAdd_6U_10U_4_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_a_int_mant_p1_2_sva,
      FpAdd_6U_10U_4_addend_larger_asn_13_mx0w1, and_dcpl_453);
  assign FpAdd_6U_10U_4_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_asn_13_mx0w1,
      FpAdd_6U_10U_4_a_int_mant_p1_2_sva, and_dcpl_453);
  assign FpAdd_6U_10U_4_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_a_int_mant_p1_3_sva,
      FpAdd_6U_10U_4_addend_larger_asn_7_mx0w1, and_dcpl_457);
  assign FpAdd_6U_10U_4_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_asn_7_mx0w1,
      FpAdd_6U_10U_4_a_int_mant_p1_3_sva, and_dcpl_457);
  assign FpAdd_6U_10U_4_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_a_int_mant_p1_sva,
      FpAdd_6U_10U_4_addend_larger_asn_1_mx0w1, and_dcpl_461);
  assign FpAdd_6U_10U_4_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_asn_1_mx0w1,
      FpAdd_6U_10U_4_a_int_mant_p1_sva, and_dcpl_461);
  assign nl_FpAdd_6U_10U_5_b_right_shift_qr_1_sva = ({reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_b_right_shift_qr_1_sva = nl_FpAdd_6U_10U_5_b_right_shift_qr_1_sva[5:0];
  assign nl_FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1 = ({reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1 = nl_FpAdd_6U_10U_5_a_right_shift_qr_1_sva_1[5:0];
  assign FpAdd_6U_10U_5_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_a_int_mant_p1_1_sva,
      FpAdd_6U_10U_5_addend_larger_asn_19_mx0w1, and_dcpl_465);
  assign FpAdd_6U_10U_5_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_asn_19_mx0w1,
      FpAdd_6U_10U_5_a_int_mant_p1_1_sva, and_dcpl_465);
  assign nl_FpAdd_6U_10U_5_b_right_shift_qr_2_sva = ({reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_b_right_shift_qr_2_sva = nl_FpAdd_6U_10U_5_b_right_shift_qr_2_sva[5:0];
  assign nl_FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1 = ({reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1 = nl_FpAdd_6U_10U_5_a_right_shift_qr_2_sva_1[5:0];
  assign FpAdd_6U_10U_5_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_a_int_mant_p1_2_sva,
      FpAdd_6U_10U_5_addend_larger_asn_13_mx0w1, and_dcpl_469);
  assign FpAdd_6U_10U_5_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_asn_13_mx0w1,
      FpAdd_6U_10U_5_a_int_mant_p1_2_sva, and_dcpl_469);
  assign nl_FpAdd_6U_10U_5_b_right_shift_qr_3_sva = ({reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_b_right_shift_qr_3_sva = nl_FpAdd_6U_10U_5_b_right_shift_qr_3_sva[5:0];
  assign nl_FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1 = ({reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1 = nl_FpAdd_6U_10U_5_a_right_shift_qr_3_sva_1[5:0];
  assign FpAdd_6U_10U_5_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_a_int_mant_p1_3_sva,
      FpAdd_6U_10U_5_addend_larger_asn_7_mx0w1, and_dcpl_473);
  assign FpAdd_6U_10U_5_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_asn_7_mx0w1,
      FpAdd_6U_10U_5_a_int_mant_p1_3_sva, and_dcpl_473);
  assign nl_FpAdd_6U_10U_5_b_right_shift_qr_sva = ({reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_b_right_shift_qr_sva = nl_FpAdd_6U_10U_5_b_right_shift_qr_sva[5:0];
  assign nl_FpAdd_6U_10U_5_a_right_shift_qr_sva_1 = ({reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp
      , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 , reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2})
      + ({(~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp) , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1)
      , (~ reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2)}) + 6'b1;
  assign FpAdd_6U_10U_5_a_right_shift_qr_sva_1 = nl_FpAdd_6U_10U_5_a_right_shift_qr_sva_1[5:0];
  assign FpAdd_6U_10U_5_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_a_int_mant_p1_sva,
      FpAdd_6U_10U_5_addend_larger_asn_1_mx0w1, and_dcpl_477);
  assign FpAdd_6U_10U_5_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_asn_1_mx0w1,
      FpAdd_6U_10U_5_a_int_mant_p1_sva, and_dcpl_477);
  assign FpAdd_6U_10U_6_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_a_int_mant_p1_1_sva,
      FpAdd_6U_10U_6_addend_larger_asn_19_mx0w1, and_dcpl_481);
  assign FpAdd_6U_10U_6_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_asn_19_mx0w1,
      FpAdd_6U_10U_6_a_int_mant_p1_1_sva, and_dcpl_481);
  assign FpAdd_6U_10U_6_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_a_int_mant_p1_2_sva,
      FpAdd_6U_10U_6_addend_larger_asn_13_mx0w1, and_dcpl_485);
  assign FpAdd_6U_10U_6_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_asn_13_mx0w1,
      FpAdd_6U_10U_6_a_int_mant_p1_2_sva, and_dcpl_485);
  assign FpAdd_6U_10U_6_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_a_int_mant_p1_3_sva,
      FpAdd_6U_10U_6_addend_larger_asn_7_mx0w1, and_dcpl_489);
  assign FpAdd_6U_10U_6_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_asn_7_mx0w1,
      FpAdd_6U_10U_6_a_int_mant_p1_3_sva, and_dcpl_489);
  assign FpAdd_6U_10U_6_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_a_int_mant_p1_sva,
      FpAdd_6U_10U_6_addend_larger_asn_1_mx0w1, and_dcpl_493);
  assign FpAdd_6U_10U_6_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_asn_1_mx0w1,
      FpAdd_6U_10U_6_a_int_mant_p1_sva, and_dcpl_493);
  assign FpAdd_6U_10U_7_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_a_int_mant_p1_1_sva,
      FpAdd_6U_10U_7_addend_larger_asn_19_mx0w1, and_dcpl_497);
  assign FpAdd_6U_10U_7_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_asn_19_mx0w1,
      FpAdd_6U_10U_7_a_int_mant_p1_1_sva, and_dcpl_497);
  assign FpAdd_6U_10U_7_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_a_int_mant_p1_2_sva,
      FpAdd_6U_10U_7_addend_larger_asn_13_mx0w1, and_dcpl_501);
  assign FpAdd_6U_10U_7_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_asn_13_mx0w1,
      FpAdd_6U_10U_7_a_int_mant_p1_2_sva, and_dcpl_501);
  assign FpAdd_6U_10U_7_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_a_int_mant_p1_3_sva,
      FpAdd_6U_10U_7_addend_larger_asn_7_mx0w1, and_dcpl_505);
  assign FpAdd_6U_10U_7_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_asn_7_mx0w1,
      FpAdd_6U_10U_7_a_int_mant_p1_3_sva, and_dcpl_505);
  assign FpAdd_6U_10U_7_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_a_int_mant_p1_sva,
      FpAdd_6U_10U_7_addend_larger_asn_1_mx0w1, and_dcpl_509);
  assign FpAdd_6U_10U_7_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_asn_1_mx0w1,
      FpAdd_6U_10U_7_a_int_mant_p1_sva, and_dcpl_509);
  assign FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_nl = FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm
      | (~ o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_nl), o_col0_1_FpMantRNE_23U_11U_4_else_and_tmp);
  assign FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_1_nl = FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm
      | (~ o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_1_nl), o_col0_2_FpMantRNE_23U_11U_4_else_and_tmp);
  assign FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_2_nl = FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm
      | (~ o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_2_nl), o_col0_3_FpMantRNE_23U_11U_4_else_and_tmp);
  assign FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_3_nl = FpAdd_6U_10U_4_is_inf_lpi_1_dfm
      | (~ o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_4_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_4_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_4_if_4_FpAdd_6U_10U_4_if_4_or_3_nl), o_col0_4_FpMantRNE_23U_11U_4_else_and_tmp);
  assign FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_nl = FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm
      | (~ o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_nl), o_col1_1_FpMantRNE_23U_11U_5_else_and_tmp);
  assign FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_1_nl = FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm
      | (~ o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_1_nl), o_col1_2_FpMantRNE_23U_11U_5_else_and_tmp);
  assign FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_2_nl = FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm
      | (~ o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_2_nl), o_col1_3_FpMantRNE_23U_11U_5_else_and_tmp);
  assign FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_3_nl = FpAdd_6U_10U_5_is_inf_lpi_1_dfm
      | (~ o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_5_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_5_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_5_if_4_FpAdd_6U_10U_5_if_4_or_3_nl), o_col1_4_FpMantRNE_23U_11U_5_else_and_tmp);
  assign FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_nl = FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm
      | (~ o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_nl), o_col2_1_FpMantRNE_23U_11U_6_else_and_tmp);
  assign FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_1_nl = FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm
      | (~ o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_1_nl), o_col2_2_FpMantRNE_23U_11U_6_else_and_tmp);
  assign FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_2_nl = FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm
      | (~ o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_2_nl), o_col2_3_FpMantRNE_23U_11U_6_else_and_tmp);
  assign FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_3_nl = FpAdd_6U_10U_6_is_inf_lpi_1_dfm
      | (~ o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_6_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_6_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_6_if_4_FpAdd_6U_10U_6_if_4_or_3_nl), o_col2_4_FpMantRNE_23U_11U_6_else_and_tmp);
  assign FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_nl = FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm
      | (~ o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm,
      (FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_nl), o_col3_1_FpMantRNE_23U_11U_7_else_and_tmp);
  assign FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_1_nl = FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm
      | (~ o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm,
      (FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_1_nl), o_col3_2_FpMantRNE_23U_11U_7_else_and_tmp);
  assign FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_2_nl = FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm
      | (~ o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm,
      (FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_2_nl), o_col3_3_FpMantRNE_23U_11U_7_else_and_tmp);
  assign FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_3_nl = FpAdd_6U_10U_7_is_inf_lpi_1_dfm
      | (~ o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_7_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_7_is_inf_lpi_1_dfm,
      (FpAdd_6U_10U_7_if_4_FpAdd_6U_10U_7_if_4_or_3_nl), o_col3_4_FpMantRNE_23U_11U_7_else_and_tmp);
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_11_m1c = ~(IsNaN_6U_10U_15_land_lpi_1_dfm_5
      | IsNaN_6U_10U_14_land_lpi_1_dfm_5);
  assign FpAdd_6U_10U_7_and_3_tmp = o_col3_4_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1
      & o_col3_4_FpMantRNE_23U_11U_7_else_and_tmp;
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_9_m1c = ~(IsNaN_6U_10U_15_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_7_and_2_tmp = o_col3_3_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1
      & o_col3_3_FpMantRNE_23U_11U_7_else_and_tmp;
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_7_m1c = ~(IsNaN_6U_10U_15_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_14_land_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_7_and_1_tmp = o_col3_2_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1
      & o_col3_2_FpMantRNE_23U_11U_7_else_and_tmp;
  assign FpAdd_6U_10U_7_FpAdd_6U_10U_7_nor_5_m1c = ~(IsNaN_6U_10U_15_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_14_land_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_7_and_tmp = o_col3_1_FpAdd_6U_10U_7_if_4_if_acc_1_itm_5_1 &
      o_col3_1_FpMantRNE_23U_11U_7_else_and_tmp;
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_11_m1c = ~(IsNaN_6U_10U_13_land_lpi_1_dfm_5
      | IsNaN_6U_10U_11_land_lpi_1_dfm_5);
  assign FpAdd_6U_10U_6_and_3_tmp = o_col2_4_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1
      & o_col2_4_FpMantRNE_23U_11U_6_else_and_tmp;
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_9_m1c = ~(IsNaN_6U_10U_13_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_11_land_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_6_and_2_tmp = o_col2_3_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1
      & o_col2_3_FpMantRNE_23U_11U_6_else_and_tmp;
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_7_m1c = ~(IsNaN_6U_10U_13_land_2_lpi_1_dfm_3
      | IsNaN_6U_10U_11_land_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_6_and_1_tmp = o_col2_2_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1
      & o_col2_2_FpMantRNE_23U_11U_6_else_and_tmp;
  assign FpAdd_6U_10U_6_FpAdd_6U_10U_6_nor_5_m1c = ~(IsNaN_6U_10U_13_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_9_land_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_6_and_tmp = o_col2_1_FpAdd_6U_10U_6_if_4_if_acc_1_itm_5_1 &
      o_col2_1_FpMantRNE_23U_11U_6_else_and_tmp;
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_11_m1c = ~(IsNaN_6U_10U_11_land_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_lpi_1_dfm_5);
  assign FpAdd_6U_10U_5_and_3_tmp = o_col1_4_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1
      & o_col1_4_FpMantRNE_23U_11U_5_else_and_tmp;
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_9_m1c = ~(IsNaN_6U_10U_11_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_5_and_2_tmp = o_col1_3_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1
      & o_col1_3_FpMantRNE_23U_11U_5_else_and_tmp;
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_7_m1c = ~(IsNaN_6U_10U_11_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_5_and_1_tmp = o_col1_2_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1
      & o_col1_2_FpMantRNE_23U_11U_5_else_and_tmp;
  assign FpAdd_6U_10U_5_FpAdd_6U_10U_5_nor_5_m1c = ~(IsNaN_6U_10U_9_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_5_and_tmp = o_col1_1_FpAdd_6U_10U_5_if_4_if_acc_1_itm_5_1 &
      o_col1_1_FpMantRNE_23U_11U_5_else_and_tmp;
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_11_m1c = ~(IsNaN_6U_10U_9_land_lpi_1_dfm_3
      | IsNaN_6U_10U_8_land_lpi_1_dfm_5);
  assign FpAdd_6U_10U_4_and_3_tmp = o_col0_4_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1
      & o_col0_4_FpMantRNE_23U_11U_4_else_and_tmp;
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_9_m1c = ~(IsNaN_6U_10U_9_land_3_lpi_1_dfm_3
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_4_and_2_tmp = o_col0_3_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1
      & o_col0_3_FpMantRNE_23U_11U_4_else_and_tmp;
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_7_m1c = ~(IsNaN_6U_10U_9_land_2_lpi_1_dfm_3
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_4_and_1_tmp = o_col0_2_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1
      & o_col0_2_FpMantRNE_23U_11U_4_else_and_tmp;
  assign FpAdd_6U_10U_4_FpAdd_6U_10U_4_nor_5_m1c = ~(IsNaN_6U_10U_9_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_4_and_tmp = o_col0_1_FpAdd_6U_10U_4_if_4_if_acc_1_itm_5_1 &
      o_col0_1_FpMantRNE_23U_11U_4_else_and_tmp;
  assign FpAdd_6U_10U_4_is_inf_1_lpi_1_dfm = ~(o_col0_1_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_4_int_mant_p1_1_sva_3[23])));
  assign FpAdd_6U_10U_4_is_inf_2_lpi_1_dfm = ~(o_col0_2_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_4_int_mant_p1_2_sva_3[23])));
  assign FpAdd_6U_10U_4_is_inf_3_lpi_1_dfm = ~(o_col0_3_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_4_int_mant_p1_3_sva_3[23])));
  assign FpAdd_6U_10U_4_is_inf_lpi_1_dfm = ~(o_col0_4_FpAdd_6U_10U_4_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_4_int_mant_p1_sva_3[23])));
  assign FpAdd_6U_10U_5_is_inf_1_lpi_1_dfm = ~(o_col1_1_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_5_int_mant_p1_1_sva_3[23])));
  assign FpAdd_6U_10U_5_is_inf_2_lpi_1_dfm = ~(o_col1_2_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_5_int_mant_p1_2_sva_3[23])));
  assign FpAdd_6U_10U_5_is_inf_3_lpi_1_dfm = ~(o_col1_3_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_5_int_mant_p1_3_sva_3[23])));
  assign FpAdd_6U_10U_5_is_inf_lpi_1_dfm = ~(o_col1_4_FpAdd_6U_10U_5_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_5_int_mant_p1_sva_3[23])));
  assign FpAdd_6U_10U_6_is_inf_1_lpi_1_dfm = ~(o_col2_1_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_6_int_mant_p1_1_sva_3[23])));
  assign FpAdd_6U_10U_6_is_inf_2_lpi_1_dfm = ~(o_col2_2_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_6_int_mant_p1_2_sva_3[23])));
  assign FpAdd_6U_10U_6_is_inf_3_lpi_1_dfm = ~(o_col2_3_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_6_int_mant_p1_3_sva_3[23])));
  assign FpAdd_6U_10U_6_is_inf_lpi_1_dfm = ~(o_col2_4_FpAdd_6U_10U_6_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_6_int_mant_p1_sva_3[23])));
  assign FpAdd_6U_10U_7_is_inf_1_lpi_1_dfm = ~(o_col3_1_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_7_int_mant_p1_1_sva_3[23])));
  assign FpAdd_6U_10U_7_is_inf_2_lpi_1_dfm = ~(o_col3_2_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_7_int_mant_p1_2_sva_3[23])));
  assign FpAdd_6U_10U_7_is_inf_3_lpi_1_dfm = ~(o_col3_3_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_7_int_mant_p1_3_sva_3[23])));
  assign FpAdd_6U_10U_7_is_inf_lpi_1_dfm = ~(o_col3_4_FpAdd_6U_10U_7_if_3_if_acc_1_itm_5_1
      | (~ (FpAdd_6U_10U_7_int_mant_p1_sva_3[23])));
  assign FpAdd_6U_10U_o_sign_or_9_nl = and_dcpl_1151 | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp)
      & and_dcpl_1153);
  assign FpAdd_6U_10U_o_sign_2_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[31]),
      (~ (chn_data_in_rsci_d_mxwt[159])), FpAdd_6U_10U_o_sign_or_9_nl);
  assign FpAdd_6U_10U_o_sign_or_6_nl = and_dcpl_1171 | ((~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp)
      & and_dcpl_1173);
  assign FpAdd_6U_10U_o_sign_3_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[47]),
      (~ (chn_data_in_rsci_d_mxwt[175])), FpAdd_6U_10U_o_sign_or_6_nl);
  assign FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_1_mx0 = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[95]),
      (chn_data_in_rsci_d_mxwt[159]), FpAdd_6U_10U_1_mux_19_mx0w2, {IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp
      , and_dcpl_1156 , and_dcpl_1158});
  assign FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_1_mx0 = MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[111]),
      (chn_data_in_rsci_d_mxwt[175]), FpAdd_6U_10U_1_mux_36_mx0w2, {IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp
      , and_dcpl_1176 , and_dcpl_1178});
  assign m_row1_if_d2_or_9_nl = and_dcpl_1161 | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp)
      & and_dcpl_1163);
  assign FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[159]),
      (~ (chn_data_in_rsci_d_mxwt[95])), m_row1_if_d2_or_9_nl);
  assign m_row1_if_d2_or_6_nl = and_dcpl_1181 | ((~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp)
      & and_dcpl_1183);
  assign FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[175]),
      (~ (chn_data_in_rsci_d_mxwt[111])), m_row1_if_d2_or_6_nl);
  assign FpAdd_6U_10U_1_o_sign_or_15_nl = and_dcpl_1166 | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp)
      & and_dcpl_1168);
  assign FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[95]),
      (~ (chn_data_in_rsci_d_mxwt[223])), FpAdd_6U_10U_1_o_sign_or_15_nl);
  assign FpAdd_6U_10U_1_o_sign_or_12_nl = and_dcpl_1186 | ((~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp)
      & and_dcpl_1188);
  assign FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[111]),
      (~ (chn_data_in_rsci_d_mxwt[239])), FpAdd_6U_10U_1_o_sign_or_12_nl);
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva = ~((z_out[17]) | (~((z_out[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva = (z_out[17]) & (~((z_out[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva = ~((z_out_15[17])
      | (~((z_out_15[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva = (z_out_15[17]) &
      (~((z_out_15[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva = ~((z_out_14[17])
      | (~((z_out_14[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva = (z_out_14[17]) &
      (~((z_out_14[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva = ~((z_out_13[17])
      | (~((z_out_13[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva = (z_out_13[17]) &
      (~((z_out_13[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva = ~((z_out_12[17])
      | (~((z_out_12[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva = (z_out_12[17]) &
      (~((z_out_12[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva = ~((z_out_11[17])
      | (~((z_out_11[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva = (z_out_11[17]) &
      (~((z_out_11[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva = ~((z_out_10[17])
      | (~((z_out_10[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva = (z_out_10[17]) &
      (~((z_out_10[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva = ~((z_out_9[17]) |
      (~((z_out_9[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva = (z_out_9[17]) & (~((z_out_9[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva = ~((z_out_8[17]) |
      (~((z_out_8[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva = (z_out_8[17]) & (~((z_out_8[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva = ~((z_out_7[17]) |
      (~((z_out_7[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva = (z_out_7[17]) & (~((z_out_7[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva = ~((z_out_6[17]) |
      (~((z_out_6[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva = (z_out_6[17]) & (~((z_out_6[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva = ~((z_out_5[17]) |
      (~((z_out_5[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva = (z_out_5[17]) & (~((z_out_5[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva = ~((z_out_4[17]) |
      (~((z_out_4[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva = (z_out_4[17]) & (~((z_out_4[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva = ~((z_out_3[17]) |
      (~((z_out_3[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva = (z_out_3[17]) & (~((z_out_3[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva = ~((z_out_2[17]) |
      (~((z_out_2[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva = (z_out_2[17]) & (~((z_out_2[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva = ~((z_out_1[17]) |
      (~((z_out_1[16:15]!=2'b00))));
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva = (z_out_1[17]) & (~((z_out_1[16:15]==2'b11)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_sva = ~((z_out[17]) | (~((z_out[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_sva = (z_out[17]) & (~((z_out[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_15_sva = ~((z_out_1[17]) |
      (~((z_out_1[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_15_sva = (z_out_1[17]) & (~((z_out_1[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_14_sva = ~((z_out_2[17]) |
      (~((z_out_2[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_14_sva = (z_out_2[17]) & (~((z_out_2[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_13_sva = ~((z_out_3[17]) |
      (~((z_out_3[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_13_sva = (z_out_3[17]) & (~((z_out_3[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_12_sva = ~((z_out_4[17]) |
      (~((z_out_4[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_12_sva = (z_out_4[17]) & (~((z_out_4[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_11_sva = ~((z_out_5[17]) |
      (~((z_out_5[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_11_sva = (z_out_5[17]) & (~((z_out_5[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_10_sva = ~((z_out_6[17]) |
      (~((z_out_6[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_10_sva = (z_out_6[17]) & (~((z_out_6[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_9_sva = ~((z_out_7[17]) | (~((z_out_7[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_9_sva = (z_out_7[17]) & (~((z_out_7[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_8_sva = ~((z_out_8[17]) | (~((z_out_8[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_8_sva = (z_out_8[17]) & (~((z_out_8[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_7_sva = ~((z_out_9[17]) | (~((z_out_9[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_7_sva = (z_out_9[17]) & (~((z_out_9[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_6_sva = ~((z_out_10[17]) |
      (~((z_out_10[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_6_sva = (z_out_10[17]) & (~((z_out_10[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_5_sva = ~((z_out_11[17]) |
      (~((z_out_11[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_5_sva = (z_out_11[17]) & (~((z_out_11[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_4_sva = ~((z_out_12[17]) |
      (~((z_out_12[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_4_sva = (z_out_12[17]) & (~((z_out_12[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_3_sva = ~((z_out_13[17]) |
      (~((z_out_13[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_3_sva = (z_out_13[17]) & (~((z_out_13[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_2_sva = ~((z_out_14[17]) |
      (~((z_out_14[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_2_sva = (z_out_14[17]) & (~((z_out_14[16:7]==10'b1111111111)));
  assign IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_1_sva = ~((z_out_15[17]) |
      (~((z_out_15[16:7]!=10'b0000000000))));
  assign IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_1_sva = (z_out_15[17]) & (~((z_out_15[16:7]==10'b1111111111)));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_nl
      = ~((chn_data_in_rsci_d_mxwt[142]) | IsZero_5U_10U_1_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_19 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_1_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_nl
      = ~((chn_data_in_rsci_d_mxwt[94]) | IsZero_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_19 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_1_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_nl
      = ~((chn_data_in_rsci_d_mxwt[158]) | IsZero_5U_10U_1_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_21 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_1_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_nl
      = ~((chn_data_in_rsci_d_mxwt[110]) | IsZero_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_21 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_nl
      = ~((chn_data_in_rsci_d_mxwt[174]) | IsZero_5U_10U_1_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_23 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_1_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_nl
      = ~((chn_data_in_rsci_d_mxwt[126]) | IsZero_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_23 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_3_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_nl
      = ~((chn_data_in_rsci_d_mxwt[190]) | IsZero_5U_10U_1_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_mux_25 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_1_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_1_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_nl
      = ~((chn_data_in_rsci_d_mxwt[78]) | IsZero_5U_10U_2_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_25 = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_2_land_1_lpi_1_dfm);
  assign m_row1_1_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2 = ~((m_row2_if_d1_mux_1_cse!=10'b0000000000));
  assign m_row1_2_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2 = ~((m_row2_if_d1_mux_4_cse!=10'b0000000000));
  assign m_row1_3_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2 = ~((m_row2_if_d1_mux_7_cse!=10'b0000000000));
  assign m_row1_4_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1!=10'b0000000000));
  assign m_row2_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign m_row2_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign m_row2_3_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign m_row2_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign IsZero_5U_10U_7_aelse_not_13 = (chn_data_in_rsci_d_mxwt[249:240]!=10'b0000000000)
      | (~ IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_sva);
  assign IsZero_5U_10U_7_aelse_not_15 = (chn_data_in_rsci_d_mxwt[233:224]!=10'b0000000000)
      | (~ IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_3_sva);
  assign IsZero_5U_10U_7_aelse_not_17 = (chn_data_in_rsci_d_mxwt[217:208]!=10'b0000000000)
      | (~ IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_2_sva);
  assign IsZero_5U_10U_7_aelse_not_19 = (chn_data_in_rsci_d_mxwt[201:192]!=10'b0000000000)
      | (~ IsZero_5U_10U_7_IsZero_5U_10U_7_nor_cse_1_sva);
  assign IsZero_5U_10U_aelse_not_13 = (chn_data_in_rsci_d_mxwt[57:48]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva);
  assign IsZero_5U_10U_aelse_not_15 = (chn_data_in_rsci_d_mxwt[41:32]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva);
  assign IsZero_5U_10U_aelse_not_17 = (chn_data_in_rsci_d_mxwt[25:16]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva);
  assign IsZero_5U_10U_aelse_not_19 = (chn_data_in_rsci_d_mxwt[9:0]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva);
  assign m_row2_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000);
  assign m_row2_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000);
  assign m_row2_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_3_mx0!=10'b0000000000);
  assign m_row2_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_2
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000);
  assign nl_m_row0_1_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_32)
      + 7'b1;
  assign m_row0_1_FpNormalize_6U_23U_acc_nl = nl_m_row0_1_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_oelse_not_9 = ((FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row0_1_FpNormalize_6U_23U_acc_nl)));
  assign nl_m_row0_2_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_33)
      + 7'b1;
  assign m_row0_2_FpNormalize_6U_23U_acc_nl = nl_m_row0_2_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_oelse_not_11 = ((FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row0_2_FpNormalize_6U_23U_acc_nl)));
  assign nl_m_row0_3_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_34)
      + 7'b1;
  assign m_row0_3_FpNormalize_6U_23U_acc_nl = nl_m_row0_3_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_oelse_not_13 = ((FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row0_3_FpNormalize_6U_23U_acc_nl)));
  assign nl_m_row0_4_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_35)
      + 7'b1;
  assign m_row0_4_FpNormalize_6U_23U_acc_nl = nl_m_row0_4_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_oelse_not_15 = ((FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row0_4_FpNormalize_6U_23U_acc_nl)));
  assign nl_m_row1_1_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_36)
      + 7'b1;
  assign m_row1_1_FpNormalize_6U_23U_1_acc_nl = nl_m_row1_1_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_9 = ((FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row1_1_FpNormalize_6U_23U_1_acc_nl)));
  assign nl_m_row1_2_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_37)
      + 7'b1;
  assign m_row1_2_FpNormalize_6U_23U_1_acc_nl = nl_m_row1_2_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_11 = ((FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row1_2_FpNormalize_6U_23U_1_acc_nl)));
  assign nl_m_row1_3_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_38)
      + 7'b1;
  assign m_row1_3_FpNormalize_6U_23U_1_acc_nl = nl_m_row1_3_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_13 = ((FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row1_3_FpNormalize_6U_23U_1_acc_nl)));
  assign nl_m_row1_4_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_39)
      + 7'b1;
  assign m_row1_4_FpNormalize_6U_23U_1_acc_nl = nl_m_row1_4_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_15 = ((FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row1_4_FpNormalize_6U_23U_1_acc_nl)));
  assign nl_m_row2_1_FpNormalize_6U_23U_2_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_40)
      + 7'b1;
  assign m_row2_1_FpNormalize_6U_23U_2_acc_nl = nl_m_row2_1_FpNormalize_6U_23U_2_acc_nl[6:0];
  assign FpNormalize_6U_23U_2_oelse_not_9 = ((FpAdd_6U_10U_2_int_mant_p1_1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row2_1_FpNormalize_6U_23U_2_acc_nl)));
  assign nl_m_row2_2_FpNormalize_6U_23U_2_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_41)
      + 7'b1;
  assign m_row2_2_FpNormalize_6U_23U_2_acc_nl = nl_m_row2_2_FpNormalize_6U_23U_2_acc_nl[6:0];
  assign FpNormalize_6U_23U_2_oelse_not_11 = ((FpAdd_6U_10U_2_int_mant_p1_2_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row2_2_FpNormalize_6U_23U_2_acc_nl)));
  assign nl_m_row2_3_FpNormalize_6U_23U_2_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_42)
      + 7'b1;
  assign m_row2_3_FpNormalize_6U_23U_2_acc_nl = nl_m_row2_3_FpNormalize_6U_23U_2_acc_nl[6:0];
  assign FpNormalize_6U_23U_2_oelse_not_13 = ((FpAdd_6U_10U_2_int_mant_p1_3_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row2_3_FpNormalize_6U_23U_2_acc_nl)));
  assign nl_m_row2_4_FpNormalize_6U_23U_2_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_43)
      + 7'b1;
  assign m_row2_4_FpNormalize_6U_23U_2_acc_nl = nl_m_row2_4_FpNormalize_6U_23U_2_acc_nl[6:0];
  assign FpNormalize_6U_23U_2_oelse_not_15 = ((FpAdd_6U_10U_2_int_mant_p1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row2_4_FpNormalize_6U_23U_2_acc_nl)));
  assign nl_m_row3_1_FpNormalize_6U_23U_3_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_44)
      + 7'b1;
  assign m_row3_1_FpNormalize_6U_23U_3_acc_nl = nl_m_row3_1_FpNormalize_6U_23U_3_acc_nl[6:0];
  assign FpNormalize_6U_23U_3_oelse_not_9 = ((FpAdd_6U_10U_3_int_mant_p1_1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row3_1_FpNormalize_6U_23U_3_acc_nl)));
  assign nl_m_row3_2_FpNormalize_6U_23U_3_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_45)
      + 7'b1;
  assign m_row3_2_FpNormalize_6U_23U_3_acc_nl = nl_m_row3_2_FpNormalize_6U_23U_3_acc_nl[6:0];
  assign FpNormalize_6U_23U_3_oelse_not_11 = ((FpAdd_6U_10U_3_int_mant_p1_2_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row3_2_FpNormalize_6U_23U_3_acc_nl)));
  assign nl_m_row3_3_FpNormalize_6U_23U_3_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_46)
      + 7'b1;
  assign m_row3_3_FpNormalize_6U_23U_3_acc_nl = nl_m_row3_3_FpNormalize_6U_23U_3_acc_nl[6:0];
  assign FpNormalize_6U_23U_3_oelse_not_13 = ((FpAdd_6U_10U_3_int_mant_p1_3_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row3_3_FpNormalize_6U_23U_3_acc_nl)));
  assign nl_m_row3_4_FpNormalize_6U_23U_3_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1) , (~ FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_47)
      + 7'b1;
  assign m_row3_4_FpNormalize_6U_23U_3_acc_nl = nl_m_row3_4_FpNormalize_6U_23U_3_acc_nl[6:0];
  assign FpNormalize_6U_23U_3_oelse_not_15 = ((FpAdd_6U_10U_3_int_mant_p1_lpi_1_dfm_mx1[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((m_row3_4_FpNormalize_6U_23U_3_acc_nl)));
  assign nl_o_col0_1_FpNormalize_6U_23U_4_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_48)
      + 7'b1;
  assign o_col0_1_FpNormalize_6U_23U_4_acc_nl = nl_o_col0_1_FpNormalize_6U_23U_4_acc_nl[6:0];
  assign FpNormalize_6U_23U_4_oelse_not_9 = ((FpAdd_6U_10U_4_int_mant_p1_1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col0_1_FpNormalize_6U_23U_4_acc_nl)));
  assign nl_o_col0_2_FpNormalize_6U_23U_4_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_49)
      + 7'b1;
  assign o_col0_2_FpNormalize_6U_23U_4_acc_nl = nl_o_col0_2_FpNormalize_6U_23U_4_acc_nl[6:0];
  assign FpNormalize_6U_23U_4_oelse_not_11 = ((FpAdd_6U_10U_4_int_mant_p1_2_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col0_2_FpNormalize_6U_23U_4_acc_nl)));
  assign nl_o_col0_3_FpNormalize_6U_23U_4_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_50)
      + 7'b1;
  assign o_col0_3_FpNormalize_6U_23U_4_acc_nl = nl_o_col0_3_FpNormalize_6U_23U_4_acc_nl[6:0];
  assign FpNormalize_6U_23U_4_oelse_not_13 = ((FpAdd_6U_10U_4_int_mant_p1_3_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col0_3_FpNormalize_6U_23U_4_acc_nl)));
  assign nl_o_col0_4_FpNormalize_6U_23U_4_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_51)
      + 7'b1;
  assign o_col0_4_FpNormalize_6U_23U_4_acc_nl = nl_o_col0_4_FpNormalize_6U_23U_4_acc_nl[6:0];
  assign FpNormalize_6U_23U_4_oelse_not_15 = ((FpAdd_6U_10U_4_int_mant_p1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col0_4_FpNormalize_6U_23U_4_acc_nl)));
  assign nl_o_col1_1_FpNormalize_6U_23U_5_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_52)
      + 7'b1;
  assign o_col1_1_FpNormalize_6U_23U_5_acc_nl = nl_o_col1_1_FpNormalize_6U_23U_5_acc_nl[6:0];
  assign FpNormalize_6U_23U_5_oelse_not_9 = ((FpAdd_6U_10U_5_int_mant_p1_1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col1_1_FpNormalize_6U_23U_5_acc_nl)));
  assign nl_o_col1_2_FpNormalize_6U_23U_5_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_53)
      + 7'b1;
  assign o_col1_2_FpNormalize_6U_23U_5_acc_nl = nl_o_col1_2_FpNormalize_6U_23U_5_acc_nl[6:0];
  assign FpNormalize_6U_23U_5_oelse_not_11 = ((FpAdd_6U_10U_5_int_mant_p1_2_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col1_2_FpNormalize_6U_23U_5_acc_nl)));
  assign nl_o_col1_3_FpNormalize_6U_23U_5_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_54)
      + 7'b1;
  assign o_col1_3_FpNormalize_6U_23U_5_acc_nl = nl_o_col1_3_FpNormalize_6U_23U_5_acc_nl[6:0];
  assign FpNormalize_6U_23U_5_oelse_not_13 = ((FpAdd_6U_10U_5_int_mant_p1_3_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col1_3_FpNormalize_6U_23U_5_acc_nl)));
  assign nl_o_col1_4_FpNormalize_6U_23U_5_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_55)
      + 7'b1;
  assign o_col1_4_FpNormalize_6U_23U_5_acc_nl = nl_o_col1_4_FpNormalize_6U_23U_5_acc_nl[6:0];
  assign FpNormalize_6U_23U_5_oelse_not_15 = ((FpAdd_6U_10U_5_int_mant_p1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col1_4_FpNormalize_6U_23U_5_acc_nl)));
  assign nl_o_col2_1_FpNormalize_6U_23U_6_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_56)
      + 7'b1;
  assign o_col2_1_FpNormalize_6U_23U_6_acc_nl = nl_o_col2_1_FpNormalize_6U_23U_6_acc_nl[6:0];
  assign FpNormalize_6U_23U_6_oelse_not_9 = ((FpAdd_6U_10U_6_int_mant_p1_1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col2_1_FpNormalize_6U_23U_6_acc_nl)));
  assign nl_o_col2_2_FpNormalize_6U_23U_6_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_57)
      + 7'b1;
  assign o_col2_2_FpNormalize_6U_23U_6_acc_nl = nl_o_col2_2_FpNormalize_6U_23U_6_acc_nl[6:0];
  assign FpNormalize_6U_23U_6_oelse_not_11 = ((FpAdd_6U_10U_6_int_mant_p1_2_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col2_2_FpNormalize_6U_23U_6_acc_nl)));
  assign nl_o_col2_3_FpNormalize_6U_23U_6_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_58)
      + 7'b1;
  assign o_col2_3_FpNormalize_6U_23U_6_acc_nl = nl_o_col2_3_FpNormalize_6U_23U_6_acc_nl[6:0];
  assign FpNormalize_6U_23U_6_oelse_not_13 = ((FpAdd_6U_10U_6_int_mant_p1_3_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col2_3_FpNormalize_6U_23U_6_acc_nl)));
  assign nl_o_col2_4_FpNormalize_6U_23U_6_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_59)
      + 7'b1;
  assign o_col2_4_FpNormalize_6U_23U_6_acc_nl = nl_o_col2_4_FpNormalize_6U_23U_6_acc_nl[6:0];
  assign FpNormalize_6U_23U_6_oelse_not_15 = ((FpAdd_6U_10U_6_int_mant_p1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col2_4_FpNormalize_6U_23U_6_acc_nl)));
  assign nl_o_col3_1_FpNormalize_6U_23U_7_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_60)
      + 7'b1;
  assign o_col3_1_FpNormalize_6U_23U_7_acc_nl = nl_o_col3_1_FpNormalize_6U_23U_7_acc_nl[6:0];
  assign FpNormalize_6U_23U_7_oelse_not_9 = ((FpAdd_6U_10U_7_int_mant_p1_1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col3_1_FpNormalize_6U_23U_7_acc_nl)));
  assign nl_o_col3_2_FpNormalize_6U_23U_7_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_61)
      + 7'b1;
  assign o_col3_2_FpNormalize_6U_23U_7_acc_nl = nl_o_col3_2_FpNormalize_6U_23U_7_acc_nl[6:0];
  assign FpNormalize_6U_23U_7_oelse_not_11 = ((FpAdd_6U_10U_7_int_mant_p1_2_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col3_2_FpNormalize_6U_23U_7_acc_nl)));
  assign nl_o_col3_3_FpNormalize_6U_23U_7_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_62)
      + 7'b1;
  assign o_col3_3_FpNormalize_6U_23U_7_acc_nl = nl_o_col3_3_FpNormalize_6U_23U_7_acc_nl[6:0];
  assign FpNormalize_6U_23U_7_oelse_not_13 = ((FpAdd_6U_10U_7_int_mant_p1_3_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col3_3_FpNormalize_6U_23U_7_acc_nl)));
  assign nl_o_col3_4_FpNormalize_6U_23U_7_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp)
      , (~ reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1) , (~ reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_8687f6a8ea077364acb8a832561c79a95444_63)
      + 7'b1;
  assign o_col3_4_FpNormalize_6U_23U_7_acc_nl = nl_o_col3_4_FpNormalize_6U_23U_7_acc_nl[6:0];
  assign FpNormalize_6U_23U_7_oelse_not_15 = ((FpAdd_6U_10U_7_int_mant_p1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((o_col3_4_FpNormalize_6U_23U_7_acc_nl)));
  assign m_row0_asn_184 = IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_186 = IsNaN_6U_10U_14_land_2_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_188 = IsNaN_6U_10U_14_land_1_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_190 = IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_192 = IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_194 = IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_196 = IsNaN_6U_10U_10_land_3_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_198 = IsNaN_6U_10U_10_land_2_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_200 = IsNaN_6U_10U_10_land_1_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_202 = IsNaN_6U_10U_8_land_3_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_204 = IsNaN_6U_10U_8_land_2_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_206 = IsNaN_6U_10U_8_land_1_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_208 = IsNaN_6U_10U_14_land_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_210 = IsNaN_6U_10U_11_land_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_212 = IsNaN_6U_10U_10_land_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_asn_214 = IsNaN_6U_10U_8_land_lpi_1_dfm_5 & (~ m_row0_unequal_tmp_4);
  assign m_row0_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      = (m_row2_if_d1_mux_1_cse!=10'b0000000000);
  assign m_row0_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      = (m_row2_if_d1_mux_4_cse!=10'b0000000000);
  assign m_row0_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      = (m_row2_if_d1_mux_7_cse!=10'b0000000000);
  assign m_row0_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_2
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_3_mx1!=10'b0000000000);
  assign and_dcpl_3 = (cfg_precision[1]) & main_stage_v_4 & or_181_cse;
  assign and_dcpl_52 = or_181_cse & (cfg_precision==2'b10) & chn_data_in_rsci_bawt;
  assign or_dcpl_1 = (cfg_precision!=2'b10);
  assign and_dcpl_57 = reg_chn_data_out_rsci_ld_core_psct_cse & chn_data_in_rsci_bawt;
  assign not_tmp_35 = ~(nor_562_cse | (cfg_precision!=2'b10));
  assign or_tmp_5 = IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign or_tmp_8 = IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp;
  assign nand_tmp_2 = ~(chn_data_in_rsci_bawt & not_tmp_35);
  assign and_72_cse = IsNaN_6U_10U_land_2_lpi_1_dfm & or_dcpl_1;
  assign or_tmp_16 = IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
  assign or_tmp_19 = IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp | IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign or_tmp_22 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign or_tmp_25 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign nand_tmp_15 = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign or_tmp_27 = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign nand_tmp_16 = ~(or_tmp_27 & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_tmp_30 = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign or_tmp_33 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign or_tmp_36 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign or_tmp_39 = IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign or_tmp_42 = IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign nand_tmp_31 = ~((~(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign or_tmp_44 = IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign or_tmp_45 = IsNaN_6U_10U_6_land_1_lpi_1_dfm | and_dcpl_52;
  assign and_tmp_1 = IsNaN_6U_10U_6_land_1_lpi_1_dfm & nand_tmp_2;
  assign mux_tmp_35 = MUX_s_1_2_2(and_tmp_1, or_tmp_45, or_tmp_44);
  assign or_tmp_48 = IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign or_tmp_52 = IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign or_tmp_57 = IsNaN_6U_10U_7_land_3_lpi_1_dfm | IsNaN_6U_10U_6_land_3_lpi_1_dfm;
  assign or_tmp_65 = IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign or_87_cse = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | main_stage_v_1;
  assign mux_tmp_49 = MUX_s_1_2_2(nor_546_cse, or_87_cse, chn_data_in_rsci_bawt);
  assign nor_559_cse = ~((~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_3) | reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse);
  assign or_92_nl = nor_559_cse | reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse;
  assign mux_tmp_51 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_92_nl);
  assign not_tmp_81 = ~((~(nor_559_cse | reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_555_cse = ~((~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_3) | reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse);
  assign or_102_nl = nor_555_cse | reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse;
  assign mux_tmp_56 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_102_nl);
  assign not_tmp_83 = ~((~(nor_555_cse | reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_551_cse = ~((~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_3) | reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse);
  assign or_112_nl = nor_551_cse | reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse;
  assign mux_tmp_61 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_112_nl);
  assign not_tmp_85 = ~((~(nor_551_cse | reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_545_cse = ~((~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_3) | reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse);
  assign or_127_nl = nor_545_cse | reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse;
  assign mux_tmp_69 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_127_nl);
  assign not_tmp_90 = ~((~(nor_545_cse | reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_tmp_72 = FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_2_cse & main_stage_v_1;
  assign mux_tmp_73 = MUX_s_1_2_2(nor_tmp_72, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_92 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_72));
  assign mux_74_nl = MUX_s_1_2_2(not_tmp_92, mux_tmp_73, or_tmp_52);
  assign mux_75_nl = MUX_s_1_2_2(not_tmp_92, mux_tmp_73, or_tmp_57);
  assign mux_tmp_76 = MUX_s_1_2_2((mux_75_nl), (mux_74_nl), nor_57_cse);
  assign nor_540_cse = ~((~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_3) | reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse);
  assign or_145_nl = nor_540_cse | reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse;
  assign mux_tmp_81 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_145_nl);
  assign not_tmp_96 = ~((~(nor_540_cse | reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_tmp_78 = FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_3_cse & main_stage_v_1;
  assign mux_tmp_85 = MUX_s_1_2_2(nor_tmp_78, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_98 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_78));
  assign mux_86_nl = MUX_s_1_2_2(not_tmp_98, mux_tmp_85, or_tmp_48);
  assign mux_87_nl = MUX_s_1_2_2(not_tmp_98, mux_tmp_85, or_152_cse);
  assign mux_tmp_88 = MUX_s_1_2_2((mux_87_nl), (mux_86_nl), nor_57_cse);
  assign nor_535_cse = ~((~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_3) | reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse);
  assign or_163_nl = nor_535_cse | reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse;
  assign mux_tmp_93 = MUX_s_1_2_2(main_stage_en_1, mux_79_cse, or_163_nl);
  assign not_tmp_102 = ~((~(nor_535_cse | reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse))
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_1));
  assign nor_tmp_84 = FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_4_cse & main_stage_v_1;
  assign mux_tmp_97 = MUX_s_1_2_2(nor_tmp_84, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_104 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_84));
  assign mux_98_nl = MUX_s_1_2_2(not_tmp_104, mux_tmp_97, or_tmp_44);
  assign or_176_nl = IsNaN_6U_10U_6_land_1_lpi_1_dfm | IsNaN_6U_10U_7_land_1_lpi_1_dfm;
  assign mux_99_nl = MUX_s_1_2_2(not_tmp_104, mux_tmp_97, or_176_nl);
  assign mux_tmp_100 = MUX_s_1_2_2((mux_99_nl), (mux_98_nl), nor_57_cse);
  assign or_tmp_170 = and_2591_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_109 = or_1963_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign or_tmp_183 = and_2588_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_112 = or_1962_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign or_tmp_196 = and_2585_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_115 = or_1961_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign or_tmp_211 = and_2582_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_120 = or_1960_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign mux_139_nl = MUX_s_1_2_2(not_tmp_120, or_tmp_211, or_tmp_27);
  assign mux_140_nl = MUX_s_1_2_2(not_tmp_120, or_tmp_211, or_224_cse);
  assign mux_141_nl = MUX_s_1_2_2((mux_140_nl), (mux_139_nl), nor_57_cse);
  assign mux_tmp_142 = MUX_s_1_2_2(not_tmp_120, (mux_141_nl), chn_data_in_rsci_bawt);
  assign or_tmp_224 = and_2579_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_123 = or_1959_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign mux_148_nl = MUX_s_1_2_2(not_tmp_123, or_tmp_224, or_tmp_25);
  assign mux_149_nl = MUX_s_1_2_2(not_tmp_123, or_tmp_224, or_237_cse);
  assign mux_150_nl = MUX_s_1_2_2((mux_149_nl), (mux_148_nl), nor_57_cse);
  assign mux_tmp_151 = MUX_s_1_2_2(not_tmp_123, (mux_150_nl), chn_data_in_rsci_bawt);
  assign nor_tmp_118 = reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
      & main_stage_v_1;
  assign or_tmp_243 = and_2576_cse | (~ reg_chn_data_out_rsci_ld_core_psct_cse) |
      chn_data_out_rsci_bawt;
  assign not_tmp_128 = or_1958_cse & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign mux_159_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_243, or_tmp_22);
  assign mux_160_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_243, or_256_cse);
  assign mux_161_nl = MUX_s_1_2_2((mux_160_nl), (mux_159_nl), nor_57_cse);
  assign mux_tmp_162 = MUX_s_1_2_2(not_tmp_128, (mux_161_nl), chn_data_in_rsci_bawt);
  assign nor_tmp_127 = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_2_cse & main_stage_v_1;
  assign mux_tmp_169 = MUX_s_1_2_2(nor_tmp_127, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_134 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_127));
  assign mux_170_nl = MUX_s_1_2_2(not_tmp_134, mux_tmp_169, or_tmp_16);
  assign mux_171_nl = MUX_s_1_2_2(not_tmp_134, mux_tmp_169, or_119_cse);
  assign mux_tmp_172 = MUX_s_1_2_2((mux_171_nl), (mux_170_nl), nor_57_cse);
  assign nor_tmp_130 = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_3_cse & main_stage_v_1;
  assign mux_tmp_176 = MUX_s_1_2_2(nor_tmp_130, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_138 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_130));
  assign mux_177_nl = MUX_s_1_2_2(not_tmp_138, mux_tmp_176, or_tmp_8);
  assign mux_178_nl = MUX_s_1_2_2(not_tmp_138, mux_tmp_176, or_109_cse);
  assign mux_tmp_179 = MUX_s_1_2_2((mux_178_nl), (mux_177_nl), nor_57_cse);
  assign nor_tmp_133 = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_4_cse & main_stage_v_1;
  assign mux_tmp_183 = MUX_s_1_2_2(nor_tmp_133, chn_data_in_rsci_bawt, or_181_cse);
  assign not_tmp_142 = ~((~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ nor_tmp_133));
  assign mux_184_nl = MUX_s_1_2_2(not_tmp_142, mux_tmp_183, or_tmp_5);
  assign mux_185_nl = MUX_s_1_2_2(not_tmp_142, mux_tmp_183, or_99_cse);
  assign mux_tmp_186 = MUX_s_1_2_2((mux_185_nl), (mux_184_nl), nor_57_cse);
  assign mux_tmp_191 = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_181_cse);
  assign mux_tmp_192 = MUX_s_1_2_2(and_2495_cse, and_2491_cse, or_181_cse);
  assign mux_tmp_193 = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_181_cse);
  assign not_tmp_148 = ~((cfg_precision[1]) & main_stage_v_1);
  assign or_tmp_286 = (cfg_precision[0]) | not_tmp_148;
  assign mux_tmp_198 = MUX_s_1_2_2(or_tmp_286, m_row0_unequal_tmp_3, main_stage_v_2);
  assign or_tmp_287 = and_2491_cse | mux_tmp_198;
  assign or_tmp_288 = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (cfg_precision[1]);
  assign mux_tmp_200 = MUX_s_1_2_2(mux_tmp_198, or_tmp_288, and_2491_cse);
  assign mux_tmp_201 = MUX_s_1_2_2(or_796_cse, m_row0_unequal_tmp_4, main_stage_v_3);
  assign or_tmp_290 = and_2495_cse | mux_tmp_201;
  assign mux_tmp_202 = MUX_s_1_2_2(or_tmp_290, mux_tmp_200, or_181_cse);
  assign or_310_nl = m_row0_unequal_tmp_3 | (~ (cfg_precision[1]));
  assign mux_tmp_203 = MUX_s_1_2_2(or_tmp_286, (or_310_nl), main_stage_v_2);
  assign mux_tmp_204 = MUX_s_1_2_2(mux_tmp_198, mux_tmp_203, and_2491_cse);
  assign mux_tmp_205 = MUX_s_1_2_2(or_tmp_290, mux_tmp_204, or_181_cse);
  assign mux_tmp_206 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_311_cse);
  assign mux_tmp_207 = MUX_s_1_2_2(mux_tmp_201, mux_tmp_200, or_181_cse);
  assign mux_tmp_208 = MUX_s_1_2_2(mux_tmp_201, mux_tmp_204, or_181_cse);
  assign mux_tmp_212 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_315_cse);
  assign or_tmp_302 = data_truncate_nor_tmp_5 | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_303 = and_2555_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_325_cse = nor_562_cse | m_row0_unequal_tmp_3;
  assign and_2556_cse = or_181_cse & m_row0_unequal_tmp_3;
  assign or_323_nl = and_2555_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_219 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_323_nl);
  assign or_tmp_319 = data_truncate_nor_tmp_5 | data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_320 = and_2550_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_340_nl = and_2550_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_228 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_340_nl);
  assign or_tmp_336 = data_truncate_nor_tmp_5 | data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_337 = and_2545_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_357_nl = and_2545_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_237 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_357_nl);
  assign mux_tmp_246 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_371_cse);
  assign mux_tmp_250 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_373_cse);
  assign mux_tmp_254 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_375_cse);
  assign or_tmp_359 = data_truncate_nor_tmp_5 | data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_360 = and_2537_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_380_nl = and_2537_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_258 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_380_nl);
  assign or_tmp_376 = data_truncate_nor_tmp_5 | data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_377 = and_2532_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_397_nl = and_2532_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_267 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_397_nl);
  assign or_tmp_393 = data_truncate_nor_tmp_5 | data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_394 = and_2527_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_414_nl = and_2527_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_276 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_414_nl);
  assign mux_tmp_291 = MUX_s_1_2_2(mux_tmp_204, mux_tmp_200, data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_tmp_419 = data_truncate_nor_tmp_5 | data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_420 = and_2517_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_440_nl = and_2517_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_299 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_440_nl);
  assign or_tmp_437 = main_stage_v_3 | mux_tmp_198;
  assign mux_tmp_308 = MUX_s_1_2_2(mux_tmp_198, or_tmp_288, main_stage_v_3);
  assign mux_310_nl = MUX_s_1_2_2(mux_tmp_198, mux_tmp_203, main_stage_v_3);
  assign mux_tmp_311 = MUX_s_1_2_2((mux_310_nl), or_tmp_437, data_truncate_nor_tmp_4);
  assign or_454_nl = data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_309_nl = MUX_s_1_2_2(mux_tmp_308, or_tmp_437, or_454_nl);
  assign mux_312_nl = MUX_s_1_2_2(or_tmp_287, mux_tmp_311, data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st);
  assign mux_tmp_313 = MUX_s_1_2_2((mux_312_nl), (mux_309_nl), data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_tmp_438 = main_stage_v_4 | mux_tmp_201;
  assign or_tmp_441 = data_truncate_nor_tmp_5 | data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_442 = and_2512_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_462_nl = and_2512_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_317 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_462_nl);
  assign mux_tmp_329 = MUX_s_1_2_2(mux_tmp_204, mux_tmp_200, data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_tmp_465 = data_truncate_nor_tmp_5 | data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_466 = and_2503_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_486_nl = and_2503_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_340 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_486_nl);
  assign or_500_nl = data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_349_nl = MUX_s_1_2_2(mux_tmp_308, or_tmp_437, or_500_nl);
  assign mux_350_nl = MUX_s_1_2_2(or_tmp_287, mux_tmp_311, data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st);
  assign mux_tmp_351 = MUX_s_1_2_2((mux_350_nl), (mux_349_nl), data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_tmp_485 = data_truncate_nor_tmp_5 | data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_486 = and_2498_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_506_nl = and_2498_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_355 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_506_nl);
  assign and_2496_nl = m_row0_unequal_tmp_3 & main_stage_v_2;
  assign mux_tmp_364 = MUX_s_1_2_2(or_796_cse, (and_2496_nl), nor_150_cse);
  assign or_tmp_510 = IsNaN_6U_10U_16_nor_15_itm_2 | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm_2;
  assign or_tmp_513 = data_truncate_nor_tmp_5 | data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_514 = and_2487_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_534_nl = and_2487_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_371 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_534_nl);
  assign mux_tmp_380 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_548_cse);
  assign or_tmp_532 = data_truncate_nor_tmp_5 | data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_533 = and_2481_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_553_nl = and_2481_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_384 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_553_nl);
  assign mux_tmp_393 = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_567_cse);
  assign or_tmp_551 = data_truncate_nor_tmp_5 | data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_552 = and_2475_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_572_nl = and_2475_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_397 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_572_nl);
  assign or_tmp_576 = IsNaN_6U_10U_16_nor_12_itm_2 | IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm_2;
  assign or_tmp_579 = data_truncate_nor_tmp_5 | data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign or_tmp_580 = and_2464_cse | m_row0_unequal_tmp_4 | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign or_600_nl = and_2464_cse | m_row0_unequal_tmp_4;
  assign mux_tmp_413 = MUX_s_1_2_2(and_2556_cse, or_325_cse, or_600_nl);
  assign nand_tmp_61 = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp | (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp)
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign or_620_nl = (IsNaN_6U_10U_1_land_lpi_1_dfm_3 & main_stage_v_1) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign mux_tmp_429 = MUX_s_1_2_2((or_620_nl), or_87_cse, reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse);
  assign and_2636_nl = IsNaN_6U_10U_1_land_lpi_1_dfm_3 & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign not_tmp_203 = MUX_s_1_2_2((and_2636_nl), nor_546_cse, reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse);
  assign or_626_nl = (IsNaN_6U_10U_7_land_lpi_1_dfm_3 & main_stage_v_1) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt;
  assign mux_tmp_435 = MUX_s_1_2_2((or_626_nl), or_87_cse, reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse);
  assign and_2634_nl = IsNaN_6U_10U_7_land_lpi_1_dfm_3 & main_stage_v_1 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt);
  assign not_tmp_204 = MUX_s_1_2_2((and_2634_nl), nor_546_cse, reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse);
  assign or_tmp_614 = (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse & main_stage_v_1)
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt;
  assign not_tmp_205 = FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_1_cse & main_stage_v_1
      & reg_chn_data_out_rsci_ld_core_psct_cse & (~ chn_data_out_rsci_bawt);
  assign and_2457_nl = or_tmp_65 & chn_data_in_rsci_bawt;
  assign mux_441_nl = MUX_s_1_2_2(not_tmp_205, or_tmp_614, and_2457_nl);
  assign and_2458_nl = or_629_cse & chn_data_in_rsci_bawt;
  assign mux_442_nl = MUX_s_1_2_2(not_tmp_205, or_tmp_614, and_2458_nl);
  assign mux_tmp_443 = MUX_s_1_2_2((mux_442_nl), (mux_441_nl), nor_57_cse);
  assign or_tmp_624 = (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse & main_stage_v_1)
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt;
  assign not_tmp_208 = FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_1_cse & main_stage_v_1
      & reg_chn_data_out_rsci_ld_core_psct_cse & (~ chn_data_out_rsci_bawt);
  assign or_tmp_634 = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse & main_stage_v_1)
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt;
  assign not_tmp_211 = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_1_cse & main_stage_v_1
      & reg_chn_data_out_rsci_ld_core_psct_cse & (~ chn_data_out_rsci_bawt);
  assign mux_454_nl = MUX_s_1_2_2(not_tmp_211, or_tmp_634, or_tmp_30);
  assign mux_455_nl = MUX_s_1_2_2(not_tmp_211, or_tmp_634, or_648_cse);
  assign mux_456_nl = MUX_s_1_2_2((mux_455_nl), (mux_454_nl), nor_57_cse);
  assign mux_tmp_457 = MUX_s_1_2_2(not_tmp_211, (mux_456_nl), chn_data_in_rsci_bawt);
  assign or_tmp_640 = (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse & main_stage_v_1)
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt;
  assign not_tmp_212 = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_1_cse & main_stage_v_1
      & reg_chn_data_out_rsci_ld_core_psct_cse & (~ chn_data_out_rsci_bawt);
  assign and_2449_nl = or_tmp_19 & chn_data_in_rsci_bawt;
  assign mux_458_nl = MUX_s_1_2_2(not_tmp_212, or_tmp_640, and_2449_nl);
  assign and_2450_nl = or_623_cse & chn_data_in_rsci_bawt;
  assign mux_459_nl = MUX_s_1_2_2(not_tmp_212, or_tmp_640, and_2450_nl);
  assign mux_tmp_460 = MUX_s_1_2_2((mux_459_nl), (mux_458_nl), nor_57_cse);
  assign and_tmp_56 = or_181_cse & main_stage_v_1;
  assign or_tmp_721 = IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_12_land_2_lpi_1_dfm_4)
      | IsNaN_6U_10U_10_land_2_lpi_1_dfm_4;
  assign or_tmp_723 = IsNaN_6U_10U_9_nor_1_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm_2;
  assign or_tmp_736 = IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_12_land_3_lpi_1_dfm_4)
      | IsNaN_6U_10U_10_land_3_lpi_1_dfm_4;
  assign or_tmp_738 = IsNaN_6U_10U_9_nor_2_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm_2;
  assign or_tmp_751 = IsNaN_6U_10U_10_land_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_12_land_lpi_1_dfm_4)
      | IsNaN_6U_10U_10_land_lpi_1_dfm_4;
  assign or_tmp_753 = IsNaN_6U_10U_9_nor_3_itm_2 | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm_2;
  assign or_tmp_774 = IsNaN_6U_10U_10_land_2_lpi_1_dfm_4 | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st;
  assign or_tmp_823 = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ main_stage_v_3) | m_row0_unequal_tmp_4;
  assign or_843_nl = (~ main_stage_v_3) | m_row0_unequal_tmp_4;
  assign mux_tmp_570 = MUX_s_1_2_2((or_843_nl), or_796_cse, or_181_cse);
  assign or_tmp_828 = nor_562_cse | (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign mux_tmp_603 = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_286, or_181_cse);
  assign or_tmp_923 = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ main_stage_v_2);
  assign mux_tmp_622 = MUX_s_1_2_2(or_796_cse, or_tmp_286, or_181_cse);
  assign or_tmp_963 = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign or_tmp_966 = nor_562_cse | (cfg_precision[0]) | not_tmp_148;
  assign or_tmp_976 = (~ main_stage_v_2) | IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3;
  assign or_tmp_977 = (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt
      | (~ main_stage_v_2) | IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3;
  assign and_dcpl_64 = (~ chn_data_out_rsci_bawt) & reg_chn_data_out_rsci_ld_core_psct_cse;
  assign and_dcpl_66 = or_181_cse & main_stage_v_4;
  assign and_dcpl_68 = (~ main_stage_v_4) & chn_data_out_rsci_bawt & reg_chn_data_out_rsci_ld_core_psct_cse;
  assign or_dcpl_21 = (cfg_precision[0]) | (~ chn_data_in_rsci_bawt);
  assign or_dcpl_23 = and_dcpl_64 | (~ (cfg_precision[1]));
  assign and_dcpl_74 = or_181_cse & (cfg_precision[1]);
  assign and_dcpl_78 = or_dcpl_1 & or_181_cse;
  assign and_dcpl_79 = ~((cfg_precision[0]) | IsNaN_6U_10U_IsNaN_6U_10U_and_tmp);
  assign and_dcpl_81 = (chn_data_in_rsci_d_mxwt[139:138]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_86 = IsDenorm_5U_10U_1_or_tmp & (chn_data_in_rsci_d_mxwt[142:141]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[140]);
  assign and_dcpl_88 = (cfg_precision==2'b10);
  assign or_dcpl_64 = (~(IsDenorm_5U_10U_1_or_tmp & (chn_data_in_rsci_d_mxwt[142:141]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[140:138]!=3'b111);
  assign and_dcpl_90 = or_dcpl_64 & or_181_cse;
  assign and_dcpl_92 = (~ (cfg_precision[0])) & IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign and_dcpl_94 = (chn_data_in_rsci_d_mxwt[10]) & IsDenorm_5U_10U_or_tmp & (cfg_precision[1]);
  assign and_dcpl_99 = (chn_data_in_rsci_d_mxwt[14:12]==3'b111) & or_181_cse & (chn_data_in_rsci_d_mxwt[11]);
  assign and_dcpl_101 = and_dcpl_88 & IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign or_dcpl_69 = (chn_data_in_rsci_d_mxwt[14:12]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[11:10]==2'b11)
      & IsDenorm_5U_10U_or_tmp));
  assign and_dcpl_102 = or_dcpl_69 & or_181_cse;
  assign and_dcpl_104 = and_dcpl_74 & and_dcpl_79;
  assign or_dcpl_70 = or_dcpl_1 | IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign and_dcpl_110 = ~((cfg_precision[0]) | IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp);
  assign and_dcpl_112 = (chn_data_in_rsci_d_mxwt[154]) & IsDenorm_5U_10U_1_or_1_tmp
      & (cfg_precision[1]);
  assign and_dcpl_117 = (chn_data_in_rsci_d_mxwt[158:156]==3'b111) & or_181_cse &
      (chn_data_in_rsci_d_mxwt[155]);
  assign or_dcpl_75 = (chn_data_in_rsci_d_mxwt[158:156]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[155:154]==2'b11)
      & IsDenorm_5U_10U_1_or_1_tmp));
  assign and_dcpl_120 = or_dcpl_75 & or_181_cse;
  assign and_dcpl_122 = (~ (cfg_precision[0])) & IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
  assign and_dcpl_124 = (chn_data_in_rsci_d_mxwt[26]) & IsDenorm_5U_10U_or_1_tmp
      & (cfg_precision[1]);
  assign and_dcpl_129 = (chn_data_in_rsci_d_mxwt[30:28]==3'b111) & or_181_cse & (chn_data_in_rsci_d_mxwt[27]);
  assign or_dcpl_80 = (chn_data_in_rsci_d_mxwt[30:28]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[27:26]==2'b11)
      & IsDenorm_5U_10U_or_1_tmp));
  assign and_dcpl_132 = or_dcpl_80 & or_181_cse;
  assign and_dcpl_134 = and_dcpl_74 & and_dcpl_110;
  assign and_dcpl_140 = ~((cfg_precision[0]) | IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp);
  assign and_dcpl_142 = (chn_data_in_rsci_d_mxwt[171:170]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_147 = IsDenorm_5U_10U_1_or_2_tmp & (chn_data_in_rsci_d_mxwt[174:173]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[172]);
  assign or_dcpl_86 = (~(IsDenorm_5U_10U_1_or_2_tmp & (chn_data_in_rsci_d_mxwt[174:173]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[172:170]!=3'b111);
  assign and_dcpl_150 = or_dcpl_86 & or_181_cse;
  assign and_dcpl_152 = (~ (cfg_precision[0])) & IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
  assign and_dcpl_154 = (chn_data_in_rsci_d_mxwt[42]) & IsDenorm_5U_10U_or_2_tmp
      & (cfg_precision[1]);
  assign and_dcpl_159 = (chn_data_in_rsci_d_mxwt[46:44]==3'b111) & or_181_cse & (chn_data_in_rsci_d_mxwt[43]);
  assign and_dcpl_161 = and_dcpl_88 & IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
  assign or_dcpl_91 = (chn_data_in_rsci_d_mxwt[46:44]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[43:42]==2'b11)
      & IsDenorm_5U_10U_or_2_tmp));
  assign and_dcpl_162 = or_dcpl_91 & or_181_cse;
  assign and_dcpl_164 = and_dcpl_74 & and_dcpl_140;
  assign or_dcpl_92 = or_dcpl_1 | IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
  assign and_dcpl_174 = ~((cfg_precision[0]) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign and_dcpl_175 = and_dcpl_74 & and_dcpl_174;
  assign or_dcpl_93 = or_dcpl_1 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign and_dcpl_181 = ~((cfg_precision[0]) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign and_dcpl_182 = and_dcpl_74 & and_dcpl_181;
  assign or_dcpl_94 = or_dcpl_1 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign and_dcpl_188 = ~((cfg_precision[0]) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign and_dcpl_189 = and_dcpl_74 & and_dcpl_188;
  assign or_dcpl_95 = or_dcpl_1 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign and_dcpl_199 = ~((cfg_precision[0]) | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp);
  assign and_dcpl_200 = and_dcpl_74 & and_dcpl_199;
  assign and_dcpl_206 = ~((cfg_precision[0]) | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign and_dcpl_207 = and_dcpl_74 & and_dcpl_206;
  assign and_dcpl_213 = ~((cfg_precision[0]) | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp);
  assign and_dcpl_214 = and_dcpl_74 & and_dcpl_213;
  assign and_dcpl_224 = ~((cfg_precision[0]) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign and_dcpl_225 = and_dcpl_74 & and_dcpl_224;
  assign or_dcpl_99 = or_dcpl_1 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign and_dcpl_231 = ~((cfg_precision[0]) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp);
  assign and_dcpl_232 = and_dcpl_74 & and_dcpl_231;
  assign or_dcpl_100 = or_dcpl_1 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign and_dcpl_238 = ~((cfg_precision[0]) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign and_dcpl_239 = and_dcpl_74 & and_dcpl_238;
  assign and_dcpl_245 = and_dcpl_88 & or_181_cse;
  assign and_dcpl_246 = (~ (cfg_precision[0])) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign and_dcpl_248 = (chn_data_in_rsci_d_mxwt[107:106]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_253 = IsDenorm_5U_10U_2_or_2_tmp & (chn_data_in_rsci_d_mxwt[110:109]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[108]);
  assign or_dcpl_106 = (~(IsDenorm_5U_10U_2_or_2_tmp & (chn_data_in_rsci_d_mxwt[110:109]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[108:106]!=3'b111);
  assign and_dcpl_256 = or_dcpl_106 & or_181_cse;
  assign and_dcpl_259 = (chn_data_in_rsci_d_mxwt[234]) & IsDenorm_5U_10U_7_or_2_tmp
      & (cfg_precision[1]);
  assign and_dcpl_264 = (chn_data_in_rsci_d_mxwt[238:236]==3'b111) & or_181_cse &
      (chn_data_in_rsci_d_mxwt[235]);
  assign or_dcpl_111 = (chn_data_in_rsci_d_mxwt[238:236]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[235:234]==2'b11)
      & IsDenorm_5U_10U_7_or_2_tmp));
  assign and_dcpl_267 = or_dcpl_111 & or_181_cse;
  assign and_dcpl_269 = and_dcpl_74 & and_dcpl_246;
  assign and_dcpl_270 = and_dcpl_78 & IsNaN_6U_10U_6_land_3_lpi_1_dfm;
  assign nor_335_nl = ~(IsNaN_6U_10U_6_land_3_lpi_1_dfm | and_dcpl_88);
  assign nand_98_nl = ~(IsNaN_6U_10U_6_land_3_lpi_1_dfm & or_dcpl_1);
  assign mux_650_nl = MUX_s_1_2_2((nand_98_nl), (nor_335_nl), IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign and_dcpl_271 = (mux_650_nl) & or_181_cse;
  assign and_dcpl_272 = (~ (cfg_precision[0])) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign and_dcpl_274 = (chn_data_in_rsci_d_mxwt[90]) & IsDenorm_5U_10U_2_or_1_tmp
      & (cfg_precision[1]);
  assign and_dcpl_279 = (chn_data_in_rsci_d_mxwt[94:92]==3'b111) & or_181_cse & (chn_data_in_rsci_d_mxwt[91]);
  assign and_dcpl_281 = and_dcpl_88 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign or_dcpl_116 = (chn_data_in_rsci_d_mxwt[94:92]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[91:90]==2'b11)
      & IsDenorm_5U_10U_2_or_1_tmp));
  assign and_dcpl_282 = or_dcpl_116 & or_181_cse;
  assign and_dcpl_285 = (chn_data_in_rsci_d_mxwt[218]) & IsDenorm_5U_10U_7_or_1_tmp
      & (cfg_precision[1]);
  assign and_dcpl_290 = (chn_data_in_rsci_d_mxwt[222:220]==3'b111) & or_181_cse &
      (chn_data_in_rsci_d_mxwt[219]);
  assign or_dcpl_121 = (chn_data_in_rsci_d_mxwt[222:220]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[219:218]==2'b11)
      & IsDenorm_5U_10U_7_or_1_tmp));
  assign and_dcpl_293 = or_dcpl_121 & or_181_cse;
  assign and_dcpl_295 = and_dcpl_74 & and_dcpl_272;
  assign and_dcpl_296 = and_dcpl_78 & IsNaN_6U_10U_6_land_2_lpi_1_dfm;
  assign mux_651_nl = MUX_s_1_2_2(and_dcpl_281, or_dcpl_100, IsNaN_6U_10U_6_land_2_lpi_1_dfm);
  assign and_dcpl_297 = (~ (mux_651_nl)) & or_181_cse;
  assign and_dcpl_298 = (~ (cfg_precision[0])) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign and_dcpl_300 = (chn_data_in_rsci_d_mxwt[75:74]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_305 = IsDenorm_5U_10U_2_or_tmp & (chn_data_in_rsci_d_mxwt[78:77]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[76]);
  assign and_dcpl_307 = and_dcpl_88 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign or_dcpl_126 = (~(IsDenorm_5U_10U_2_or_tmp & (chn_data_in_rsci_d_mxwt[78:77]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[76:74]!=3'b111);
  assign and_dcpl_308 = or_dcpl_126 & or_181_cse;
  assign and_dcpl_311 = (chn_data_in_rsci_d_mxwt[202]) & IsDenorm_5U_10U_7_or_tmp
      & (cfg_precision[1]);
  assign and_dcpl_316 = (chn_data_in_rsci_d_mxwt[206:204]==3'b111) & or_181_cse &
      (chn_data_in_rsci_d_mxwt[203]);
  assign or_dcpl_131 = (chn_data_in_rsci_d_mxwt[206:204]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[203:202]==2'b11)
      & IsDenorm_5U_10U_7_or_tmp));
  assign and_dcpl_319 = or_dcpl_131 & or_181_cse;
  assign and_dcpl_321 = and_dcpl_74 & and_dcpl_298;
  assign and_dcpl_322 = and_dcpl_78 & IsNaN_6U_10U_6_land_1_lpi_1_dfm;
  assign mux_652_nl = MUX_s_1_2_2(and_dcpl_307, or_dcpl_99, IsNaN_6U_10U_6_land_1_lpi_1_dfm);
  assign and_dcpl_323 = (~ (mux_652_nl)) & or_181_cse;
  assign and_dcpl_324 = (~ (cfg_precision[0])) & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign and_dcpl_333 = and_dcpl_74 & and_dcpl_324;
  assign and_dcpl_334 = (~ (cfg_precision[0])) & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
  assign and_dcpl_343 = and_dcpl_74 & and_dcpl_334;
  assign and_dcpl_344 = (~ (cfg_precision[0])) & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
  assign and_dcpl_353 = and_dcpl_74 & and_dcpl_344;
  assign and_dcpl_354 = (~ (cfg_precision[0])) & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign and_dcpl_357 = and_dcpl_88 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign mux_653_nl = MUX_s_1_2_2(and_dcpl_357, or_dcpl_95, IsNaN_6U_10U_2_land_3_lpi_1_dfm);
  assign and_dcpl_363 = (mux_653_nl) & or_181_cse;
  assign and_dcpl_364 = and_dcpl_78 & (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm);
  assign and_dcpl_366 = (~ (cfg_precision[0])) & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign and_dcpl_369 = and_dcpl_88 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign mux_654_nl = MUX_s_1_2_2(and_dcpl_369, or_dcpl_94, IsNaN_6U_10U_2_land_2_lpi_1_dfm);
  assign and_dcpl_375 = (mux_654_nl) & or_181_cse;
  assign and_dcpl_376 = and_dcpl_78 & (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm);
  assign and_dcpl_378 = (~ (cfg_precision[0])) & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign and_dcpl_381 = and_dcpl_88 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign mux_655_nl = MUX_s_1_2_2(and_dcpl_381, or_dcpl_93, IsNaN_6U_10U_2_land_1_lpi_1_dfm);
  assign and_dcpl_387 = (mux_655_nl) & or_181_cse;
  assign and_dcpl_388 = and_dcpl_78 & (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm);
  assign mux_tmp_656 = MUX_s_1_2_2(and_dcpl_161, or_dcpl_92, IsNaN_6U_10U_land_3_lpi_1_dfm);
  assign and_dcpl_391 = mux_tmp_656 & or_181_cse;
  assign or_1226_nl = IsNaN_6U_10U_land_2_lpi_1_dfm | and_dcpl_88;
  assign mux_tmp_657 = MUX_s_1_2_2(and_72_cse, (or_1226_nl), IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp);
  assign and_dcpl_394 = mux_tmp_657 & or_181_cse;
  assign mux_tmp_658 = MUX_s_1_2_2(and_dcpl_101, or_dcpl_70, IsNaN_6U_10U_land_1_lpi_1_dfm);
  assign and_dcpl_397 = mux_tmp_658 & or_181_cse;
  assign or_dcpl_168 = FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_itm_10_1 | (~ o_col0_1_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp);
  assign and_dcpl_449 = or_dcpl_168 & (~ FpAdd_6U_10U_4_is_a_greater_acc_itm_6_1);
  assign or_dcpl_170 = FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_itm_10_1 | (~
      o_col0_2_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp);
  assign and_dcpl_453 = or_dcpl_170 & (~ FpAdd_6U_10U_4_is_a_greater_acc_1_itm_6_1);
  assign or_dcpl_172 = FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_itm_10_1 | (~
      o_col0_3_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp);
  assign and_dcpl_457 = or_dcpl_172 & (~ FpAdd_6U_10U_4_is_a_greater_acc_2_itm_6_1);
  assign or_dcpl_174 = (~ o_col0_4_FpAdd_6U_10U_4_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_itm_10_1;
  assign and_dcpl_461 = or_dcpl_174 & (~ FpAdd_6U_10U_4_is_a_greater_acc_3_itm_6_1);
  assign or_dcpl_176 = (~ o_col1_1_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_itm_10_1;
  assign and_dcpl_465 = or_dcpl_176 & (~ FpAdd_6U_10U_5_is_a_greater_acc_itm_6_1);
  assign or_dcpl_178 = (~ o_col1_2_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_itm_10_1;
  assign and_dcpl_469 = or_dcpl_178 & (~ FpAdd_6U_10U_5_is_a_greater_acc_1_itm_6_1);
  assign or_dcpl_180 = FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_itm_10_1 | (~
      o_col1_3_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp);
  assign and_dcpl_473 = or_dcpl_180 & (~ FpAdd_6U_10U_5_is_a_greater_acc_2_itm_6_1);
  assign or_dcpl_182 = (~ o_col1_4_FpAdd_6U_10U_5_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_itm_10_1;
  assign and_dcpl_477 = or_dcpl_182 & (~ FpAdd_6U_10U_5_is_a_greater_acc_3_itm_6_1);
  assign or_dcpl_184 = FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_itm_10_1 | (~ o_col2_1_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp);
  assign and_dcpl_481 = or_dcpl_184 & (~ FpAdd_6U_10U_6_is_a_greater_acc_itm_6_1);
  assign or_dcpl_186 = FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_itm_10_1 | (~
      o_col2_2_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp);
  assign and_dcpl_485 = or_dcpl_186 & (~ FpAdd_6U_10U_6_is_a_greater_acc_1_itm_6_1);
  assign or_dcpl_188 = (~ o_col2_3_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_itm_10_1;
  assign and_dcpl_489 = or_dcpl_188 & (~ FpAdd_6U_10U_6_is_a_greater_acc_2_itm_6_1);
  assign or_dcpl_190 = (~ o_col2_4_FpAdd_6U_10U_6_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_itm_10_1;
  assign and_dcpl_493 = or_dcpl_190 & (~ FpAdd_6U_10U_6_is_a_greater_acc_3_itm_6_1);
  assign or_dcpl_192 = FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_itm_10_1 | (~ o_col3_1_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp);
  assign and_dcpl_497 = or_dcpl_192 & (~ FpAdd_6U_10U_7_is_a_greater_acc_itm_6_1);
  assign or_dcpl_194 = FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_itm_10_1 | (~
      o_col3_2_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp);
  assign and_dcpl_501 = or_dcpl_194 & (~ FpAdd_6U_10U_7_is_a_greater_acc_1_itm_6_1);
  assign or_dcpl_196 = FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_itm_10_1 | (~
      o_col3_3_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp);
  assign and_dcpl_505 = or_dcpl_196 & (~ FpAdd_6U_10U_7_is_a_greater_acc_2_itm_6_1);
  assign or_dcpl_198 = (~ o_col3_4_FpAdd_6U_10U_7_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_itm_10_1;
  assign and_dcpl_509 = or_dcpl_198 & (~ FpAdd_6U_10U_7_is_a_greater_acc_3_itm_6_1);
  assign or_dcpl_200 = ~(main_stage_v_4 & data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_203 = ~((cfg_precision[1]) & data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_206 = ~(main_stage_v_4 & data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_209 = ~((cfg_precision[1]) & data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_212 = ~(main_stage_v_4 & data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_215 = ~((cfg_precision[1]) & data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_218 = ~(main_stage_v_4 & data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_221 = ~((cfg_precision[1]) & data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_224 = ~(main_stage_v_4 & data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_227 = ~((cfg_precision[1]) & data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_230 = ~(main_stage_v_4 & data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_233 = ~((cfg_precision[1]) & data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_236 = ~(main_stage_v_4 & data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_239 = ~((cfg_precision[1]) & data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_242 = ~(main_stage_v_4 & data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_245 = ~((cfg_precision[1]) & data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_248 = ~(main_stage_v_4 & data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_251 = ~((cfg_precision[1]) & data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_254 = ~(main_stage_v_4 & data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_257 = ~((cfg_precision[1]) & data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_260 = ~(main_stage_v_4 & data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_263 = ~((cfg_precision[1]) & data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_266 = ~(main_stage_v_4 & data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_269 = ~((cfg_precision[1]) & data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_272 = ~(main_stage_v_4 & data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_275 = ~((cfg_precision[1]) & data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_278 = ~(main_stage_v_4 & data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_281 = ~((cfg_precision[1]) & data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_284 = ~(main_stage_v_4 & data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_287 = ~((cfg_precision[1]) & data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_290 = ~(main_stage_v_4 & data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_dcpl_293 = ~((cfg_precision[1]) & data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign and_dcpl_547 = or_181_cse & (~ (cfg_precision[1]));
  assign or_dcpl_296 = and_dcpl_64 | (~ main_stage_v_3);
  assign or_dcpl_301 = (~ main_stage_v_1) | (cfg_precision!=2'b10);
  assign or_dcpl_302 = or_dcpl_301 | and_dcpl_64;
  assign and_dcpl_644 = (~ (cfg_precision[0])) & chn_data_in_rsci_bawt;
  assign and_dcpl_645 = and_dcpl_644 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_tmp);
  assign and_dcpl_651 = and_dcpl_644 & IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
  assign or_dcpl_303 = or_dcpl_23 | or_dcpl_21;
  assign and_dcpl_658 = and_dcpl_74 & and_dcpl_651;
  assign and_dcpl_659 = and_dcpl_644 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp);
  assign and_dcpl_665 = and_dcpl_644 & IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
  assign and_dcpl_672 = and_dcpl_74 & and_dcpl_665;
  assign and_dcpl_673 = and_dcpl_140 & chn_data_in_rsci_bawt;
  assign and_dcpl_679 = and_dcpl_152 & chn_data_in_rsci_bawt;
  assign and_dcpl_686 = and_dcpl_74 & and_dcpl_679;
  assign and_dcpl_687 = and_dcpl_644 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
  assign and_dcpl_693 = and_dcpl_644 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign and_dcpl_701 = and_dcpl_644 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
  assign and_dcpl_707 = and_dcpl_644 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign and_dcpl_715 = and_dcpl_644 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
  assign and_dcpl_721 = and_dcpl_644 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign and_dcpl_729 = and_dcpl_644 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
  assign and_dcpl_735 = and_dcpl_644 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp);
  assign and_dcpl_742 = and_dcpl_74 & and_dcpl_735;
  assign and_dcpl_743 = and_dcpl_644 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
  assign and_dcpl_749 = and_dcpl_644 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign and_dcpl_756 = and_dcpl_74 & and_dcpl_749;
  assign and_dcpl_757 = and_dcpl_644 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
  assign and_dcpl_763 = and_dcpl_644 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp);
  assign and_dcpl_770 = and_dcpl_74 & and_dcpl_763;
  assign and_dcpl_771 = and_dcpl_644 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign and_dcpl_777 = and_dcpl_644 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign and_dcpl_785 = and_dcpl_644 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
  assign and_dcpl_791 = and_dcpl_644 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp);
  assign and_dcpl_799 = and_dcpl_644 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign and_dcpl_805 = and_dcpl_644 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign and_dcpl_817 = and_dcpl_88 & chn_data_out_rsci_bawt;
  assign and_dcpl_823 = and_dcpl_88 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp;
  assign and_dcpl_824 = and_dcpl_88 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp);
  assign and_dcpl_833 = and_dcpl_88 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp;
  assign and_dcpl_834 = and_dcpl_88 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp);
  assign and_dcpl_843 = and_dcpl_88 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp;
  assign and_dcpl_844 = and_dcpl_88 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp);
  assign and_dcpl_853 = and_dcpl_88 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp;
  assign and_dcpl_854 = and_dcpl_88 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp);
  assign and_dcpl_863 = and_dcpl_88 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp;
  assign and_dcpl_864 = and_dcpl_88 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp);
  assign and_dcpl_873 = and_dcpl_88 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp;
  assign and_dcpl_874 = and_dcpl_88 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp);
  assign and_dcpl_883 = and_dcpl_88 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp;
  assign and_dcpl_884 = and_dcpl_88 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp);
  assign and_dcpl_893 = and_dcpl_88 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp;
  assign and_dcpl_894 = and_dcpl_88 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp);
  assign and_dcpl_903 = and_dcpl_88 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp;
  assign and_dcpl_904 = and_dcpl_88 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp);
  assign and_dcpl_913 = and_dcpl_88 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp;
  assign and_dcpl_914 = and_dcpl_88 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp);
  assign and_dcpl_923 = and_dcpl_88 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp;
  assign and_dcpl_924 = and_dcpl_88 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp);
  assign and_dcpl_933 = and_dcpl_88 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp;
  assign and_dcpl_934 = and_dcpl_88 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp);
  assign and_dcpl_943 = and_dcpl_88 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp;
  assign and_dcpl_944 = and_dcpl_88 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp);
  assign and_dcpl_953 = and_dcpl_88 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp;
  assign and_dcpl_954 = and_dcpl_88 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp);
  assign and_dcpl_963 = and_dcpl_88 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp;
  assign and_dcpl_964 = and_dcpl_88 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp);
  assign and_dcpl_973 = and_dcpl_88 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp;
  assign and_dcpl_974 = and_dcpl_88 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp);
  assign and_dcpl_975 = ~((cfg_precision[0]) | IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp);
  assign and_dcpl_977 = (chn_data_in_rsci_d_mxwt[187:186]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_982 = IsDenorm_5U_10U_1_or_3_tmp & (chn_data_in_rsci_d_mxwt[190:189]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[188]);
  assign or_dcpl_336 = (~(IsDenorm_5U_10U_1_or_3_tmp & (chn_data_in_rsci_d_mxwt[190:189]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[188:186]!=3'b111);
  assign and_dcpl_985 = or_dcpl_336 & or_181_cse;
  assign and_dcpl_987 = (~ (cfg_precision[0])) & IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign and_dcpl_989 = (chn_data_in_rsci_d_mxwt[59:58]==2'b11) & (cfg_precision[1]);
  assign and_dcpl_994 = IsDenorm_5U_10U_or_3_tmp & (chn_data_in_rsci_d_mxwt[62:61]==2'b11)
      & or_181_cse & (chn_data_in_rsci_d_mxwt[60]);
  assign and_dcpl_996 = and_dcpl_88 & IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign or_dcpl_341 = (~(IsDenorm_5U_10U_or_3_tmp & (chn_data_in_rsci_d_mxwt[62:61]==2'b11)))
      | (chn_data_in_rsci_d_mxwt[60:58]!=3'b111);
  assign and_dcpl_997 = or_dcpl_341 & or_181_cse;
  assign and_dcpl_999 = and_dcpl_74 & and_dcpl_975;
  assign or_dcpl_342 = or_dcpl_1 | IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign and_dcpl_1001 = ~((cfg_precision[0]) | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign and_dcpl_1002 = and_dcpl_74 & and_dcpl_1001;
  assign or_dcpl_343 = or_dcpl_1 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  assign and_dcpl_1004 = ~((cfg_precision[0]) | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp);
  assign and_dcpl_1005 = and_dcpl_74 & and_dcpl_1004;
  assign and_dcpl_1007 = ~((cfg_precision[0]) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp);
  assign and_dcpl_1008 = and_dcpl_74 & and_dcpl_1007;
  assign or_dcpl_345 = or_dcpl_1 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign and_dcpl_1010 = (~ (cfg_precision[0])) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign and_dcpl_1012 = (chn_data_in_rsci_d_mxwt[122]) & IsDenorm_5U_10U_2_or_3_tmp
      & (cfg_precision[1]);
  assign and_dcpl_1017 = (chn_data_in_rsci_d_mxwt[126:124]==3'b111) & or_181_cse
      & (chn_data_in_rsci_d_mxwt[123]);
  assign and_dcpl_1019 = and_dcpl_88 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign or_dcpl_350 = (chn_data_in_rsci_d_mxwt[126:124]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[123:122]==2'b11)
      & IsDenorm_5U_10U_2_or_3_tmp));
  assign and_dcpl_1020 = or_dcpl_350 & or_181_cse;
  assign and_dcpl_1023 = (chn_data_in_rsci_d_mxwt[250]) & IsDenorm_5U_10U_7_or_3_tmp
      & (cfg_precision[1]);
  assign and_dcpl_1028 = (chn_data_in_rsci_d_mxwt[254:252]==3'b111) & or_181_cse
      & (chn_data_in_rsci_d_mxwt[251]);
  assign or_dcpl_355 = (chn_data_in_rsci_d_mxwt[254:252]!=3'b111) | (~((chn_data_in_rsci_d_mxwt[251:250]==2'b11)
      & IsDenorm_5U_10U_7_or_3_tmp));
  assign and_dcpl_1031 = or_dcpl_355 & or_181_cse;
  assign and_dcpl_1033 = and_dcpl_74 & and_dcpl_1010;
  assign and_dcpl_1034 = and_dcpl_78 & IsNaN_6U_10U_6_land_lpi_1_dfm_st;
  assign mux_659_nl = MUX_s_1_2_2(and_dcpl_1019, or_dcpl_345, IsNaN_6U_10U_6_land_lpi_1_dfm_st);
  assign and_dcpl_1035 = (~ (mux_659_nl)) & or_181_cse;
  assign and_dcpl_1036 = (~ (cfg_precision[0])) & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign and_dcpl_1045 = and_dcpl_74 & and_dcpl_1036;
  assign and_dcpl_1046 = (~ (cfg_precision[0])) & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  assign and_dcpl_1049 = and_dcpl_88 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  assign mux_660_nl = MUX_s_1_2_2(and_dcpl_1049, or_dcpl_343, IsNaN_6U_10U_2_land_lpi_1_dfm_st);
  assign and_dcpl_1055 = (mux_660_nl) & or_181_cse;
  assign and_dcpl_1056 = and_dcpl_78 & (~ IsNaN_6U_10U_2_land_lpi_1_dfm_st);
  assign mux_tmp_661 = MUX_s_1_2_2(and_dcpl_996, or_dcpl_342, IsNaN_6U_10U_land_lpi_1_dfm_st);
  assign and_dcpl_1059 = mux_tmp_661 & or_181_cse;
  assign and_dcpl_1061 = and_dcpl_644 & (~ IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp);
  assign and_dcpl_1067 = and_dcpl_644 & IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
  assign and_dcpl_1074 = and_dcpl_74 & and_dcpl_1067;
  assign and_dcpl_1075 = and_dcpl_644 & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
  assign and_dcpl_1081 = and_dcpl_644 & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign and_dcpl_1089 = and_dcpl_644 & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
  assign and_dcpl_1095 = and_dcpl_644 & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp);
  assign and_dcpl_1102 = and_dcpl_74 & and_dcpl_1095;
  assign and_dcpl_1103 = and_dcpl_644 & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign and_dcpl_1109 = and_dcpl_644 & (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp);
  assign and_dcpl_1119 = main_stage_v_1 & (cfg_precision==2'b10) & or_181_cse;
  assign and_dcpl_1122 = or_dcpl_301 & main_stage_v_2 & or_181_cse & (~ m_row0_unequal_tmp_3);
  assign or_dcpl_366 = (cfg_precision!=2'b01);
  assign and_dcpl_1126 = or_dcpl_366 & or_181_cse;
  assign or_dcpl_367 = (cfg_precision!=2'b00);
  assign and_dcpl_1129 = or_dcpl_367 & or_181_cse;
  assign and_dcpl_1131 = (~ IsNaN_6U_10U_IsNaN_6U_10U_and_tmp) & IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp;
  assign and_dcpl_1133 = ~(IsNaN_6U_10U_IsNaN_6U_10U_and_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp);
  assign and_dcpl_1136 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign and_dcpl_1138 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp);
  assign and_dcpl_1141 = (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign and_dcpl_1143 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp);
  assign and_dcpl_1146 = (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp) & IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp;
  assign and_dcpl_1148 = ~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp | IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp);
  assign and_dcpl_1151 = (~ IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp) & IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp;
  assign and_dcpl_1153 = ~(IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp);
  assign and_dcpl_1156 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign and_dcpl_1158 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp);
  assign and_dcpl_1161 = IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp & (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign and_dcpl_1163 = ~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp);
  assign and_dcpl_1166 = (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp) & IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp;
  assign and_dcpl_1168 = ~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp | IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp);
  assign and_dcpl_1171 = (~ IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp) & IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp;
  assign and_dcpl_1173 = ~(IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp);
  assign and_dcpl_1176 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign and_dcpl_1178 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp);
  assign and_dcpl_1181 = (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign and_dcpl_1183 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp);
  assign and_dcpl_1186 = (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp) & IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp;
  assign and_dcpl_1188 = ~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp | IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp);
  assign and_dcpl_1191 = (~ IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp) & IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp;
  assign and_dcpl_1193 = ~(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp | IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp);
  assign and_dcpl_1196 = (~ IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp) & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
  assign and_dcpl_1198 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp);
  assign and_dcpl_1201 = IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp & (~ IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign and_dcpl_1203 = ~(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp);
  assign and_dcpl_1206 = (~ IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp) & IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp;
  assign and_dcpl_1208 = ~(IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp);
  assign or_dcpl_368 = (~ main_stage_v_1) | (cfg_precision[1]);
  assign FpAdd_6U_10U_mux_3_itm = MUX_s_1_2_2((FpAdd_6U_10U_int_mant_p1_1_sva_1[23]),
      (FpAdd_6U_10U_int_mant_p1_1_sva[23]), reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_mux_20_itm = MUX_s_1_2_2((FpAdd_6U_10U_int_mant_p1_2_sva_1[23]),
      (FpAdd_6U_10U_int_mant_p1_2_sva[23]), reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_mux_37_itm = MUX_s_1_2_2((FpAdd_6U_10U_int_mant_p1_3_sva_1[23]),
      (FpAdd_6U_10U_int_mant_p1_3_sva[23]), reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_mux_69_itm = MUX_s_1_2_2((FpAdd_6U_10U_int_mant_p1_sva_1[23]),
      (FpAdd_6U_10U_int_mant_p1_sva[23]), reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_1_mux_3_itm = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_1_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_1_sva[23]), reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_mux_20_itm = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_2_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_2_sva[23]), reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_mux_37_itm = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_3_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_3_sva[23]), reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_1_mux_73_itm = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_sva[23]), reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse);
  assign FpAdd_6U_10U_2_mux_3_itm = MUX_s_1_2_2((FpAdd_6U_10U_2_int_mant_p1_1_sva_1[23]),
      (FpAdd_6U_10U_2_int_mant_p1_1_sva[23]), reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_mux_20_itm = MUX_s_1_2_2((FpAdd_6U_10U_2_int_mant_p1_2_sva_1[23]),
      (FpAdd_6U_10U_2_int_mant_p1_2_sva[23]), reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_mux_37_itm = MUX_s_1_2_2((FpAdd_6U_10U_2_int_mant_p1_3_sva_1[23]),
      (FpAdd_6U_10U_2_int_mant_p1_3_sva[23]), reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_2_mux_73_itm = MUX_s_1_2_2((FpAdd_6U_10U_2_int_mant_p1_sva_1[23]),
      (FpAdd_6U_10U_2_int_mant_p1_sva[23]), reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_mux_3_itm = MUX_s_1_2_2((FpAdd_6U_10U_3_int_mant_p1_1_sva_1[23]),
      (FpAdd_6U_10U_3_int_mant_p1_1_sva[23]), reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_mux_20_itm = MUX_s_1_2_2((FpAdd_6U_10U_3_int_mant_p1_2_sva_1[23]),
      (FpAdd_6U_10U_3_int_mant_p1_2_sva[23]), reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_mux_37_itm = MUX_s_1_2_2((FpAdd_6U_10U_3_int_mant_p1_3_sva_1[23]),
      (FpAdd_6U_10U_3_int_mant_p1_3_sva[23]), reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign FpAdd_6U_10U_3_mux_69_itm = MUX_s_1_2_2((FpAdd_6U_10U_3_int_mant_p1_sva_1[23]),
      (FpAdd_6U_10U_3_int_mant_p1_sva[23]), reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse);
  assign or_tmp_1099 = or_181_cse & chn_data_in_rsci_bawt & (fsm_output[1]);
  assign and_1769_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp
      & (fsm_output[1]);
  assign and_1771_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp)
      & (fsm_output[1]);
  assign and_1801_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp
      & (fsm_output[1]);
  assign and_1803_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp)
      & (fsm_output[1]);
  assign and_1833_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp
      & (fsm_output[1]);
  assign and_1835_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp)
      & (fsm_output[1]);
  assign and_1865_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp
      & (fsm_output[1]);
  assign and_1867_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp)
      & (fsm_output[1]);
  assign and_1895_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp
      & (fsm_output[1]);
  assign and_1897_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp)
      & (fsm_output[1]);
  assign and_1927_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp
      & (fsm_output[1]);
  assign and_1929_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp)
      & (fsm_output[1]);
  assign and_1959_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp
      & (fsm_output[1]);
  assign and_1961_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp)
      & (fsm_output[1]);
  assign and_1991_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp
      & (fsm_output[1]);
  assign and_1993_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp)
      & (fsm_output[1]);
  assign and_2021_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp
      & (fsm_output[1]);
  assign and_2023_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp)
      & (fsm_output[1]);
  assign and_2053_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp
      & (fsm_output[1]);
  assign and_2055_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp)
      & (fsm_output[1]);
  assign and_2085_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp
      & (fsm_output[1]);
  assign and_2087_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp)
      & (fsm_output[1]);
  assign and_2117_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp
      & (fsm_output[1]);
  assign and_2119_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp)
      & (fsm_output[1]);
  assign and_2147_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp
      & (fsm_output[1]);
  assign and_2149_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp)
      & (fsm_output[1]);
  assign and_2179_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp
      & (fsm_output[1]);
  assign and_2181_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp)
      & (fsm_output[1]);
  assign and_2211_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp
      & (fsm_output[1]);
  assign and_2213_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp)
      & (fsm_output[1]);
  assign and_2243_cse = and_dcpl_74 & and_dcpl_644 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp
      & (fsm_output[1]);
  assign and_2245_cse = and_dcpl_74 & and_dcpl_644 & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp)
      & (fsm_output[1]);
  assign chn_data_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign main_stage_v_1_mx0c1 = or_181_cse & main_stage_v_1 & (~ chn_data_in_rsci_bawt);
  assign main_stage_v_2_mx0c1 = (~ main_stage_v_1) & main_stage_v_2 & or_181_cse;
  assign main_stage_v_3_mx0c1 = (~ main_stage_v_2) & main_stage_v_3 & or_181_cse;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_181_cse;
  assign FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_4_is_a_greater_acc_itm_6_1) & or_dcpl_168;
  assign FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_4_is_a_greater_acc_1_itm_6_1) & or_dcpl_170;
  assign FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_4_is_a_greater_acc_2_itm_6_1) & or_dcpl_172;
  assign FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~ FpAdd_6U_10U_4_is_a_greater_acc_3_itm_6_1)
      & or_dcpl_174;
  assign FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_5_is_a_greater_acc_itm_6_1) & or_dcpl_176;
  assign FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_5_is_a_greater_acc_1_itm_6_1) & or_dcpl_178;
  assign FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_5_is_a_greater_acc_2_itm_6_1) & or_dcpl_180;
  assign FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~ FpAdd_6U_10U_5_is_a_greater_acc_3_itm_6_1)
      & or_dcpl_182;
  assign FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_6_is_a_greater_acc_itm_6_1) & or_dcpl_184;
  assign FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_6_is_a_greater_acc_1_itm_6_1) & or_dcpl_186;
  assign FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_6_is_a_greater_acc_2_itm_6_1) & or_dcpl_188;
  assign FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~ FpAdd_6U_10U_6_is_a_greater_acc_3_itm_6_1)
      & or_dcpl_190;
  assign FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_7_is_a_greater_acc_itm_6_1) & or_dcpl_192;
  assign FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_7_is_a_greater_acc_1_itm_6_1) & or_dcpl_194;
  assign FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~
      FpAdd_6U_10U_7_is_a_greater_acc_2_itm_6_1) & or_dcpl_196;
  assign FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1 = and_dcpl_245 & main_stage_v_2 & (~ FpAdd_6U_10U_7_is_a_greater_acc_3_itm_6_1)
      & or_dcpl_198;
  assign FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx0c1 = and_tmp_56 & and_dcpl_88 & (~
      reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse);
  assign FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx0c1 = and_tmp_56 & and_dcpl_88 & (~
      IsNaN_6U_10U_4_land_lpi_1_dfm_st_2);
  assign FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx0c1 = and_tmp_56 & and_dcpl_88 & (~
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_2);
  assign FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0c1 = and_tmp_56 & and_dcpl_88 & (~ reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse);
  assign FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_mx0c1 = and_1771_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp));
  assign FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_mx0c1 = and_1803_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp));
  assign FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_mx0c1 = and_1835_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp));
  assign FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_mx0c1 = and_1867_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp));
  assign FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_mx0c1 = and_1897_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp));
  assign FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_mx0c1 = and_1929_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp));
  assign FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_mx0c1 = and_1961_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp));
  assign FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_mx0c1 = and_1993_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp));
  assign FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_mx0c1 = and_2023_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp));
  assign FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_mx0c1 = and_2055_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp));
  assign FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_mx0c1 = and_2087_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp));
  assign FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_mx0c1 = and_2119_cse | (and_dcpl_817 &
      and_dcpl_57 & (~ FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp));
  assign FpAdd_6U_10U_qr_3_0_lpi_1_dfm_mx0c1 = and_2149_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp));
  assign FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_mx0c1 = and_2181_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp));
  assign FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_mx0c1 = and_2213_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp));
  assign FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_mx0c1 = and_2245_cse | (and_dcpl_817 & and_dcpl_57
      & (~ FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp));
  assign FpAdd_6U_10U_o_sign_1_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1133;
  assign FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1138;
  assign FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1143;
  assign FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1148;
  assign FpAdd_6U_10U_3_o_sign_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1193;
  assign FpAdd_6U_10U_2_o_sign_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1198;
  assign FpAdd_6U_10U_1_o_sign_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1203;
  assign FpAdd_6U_10U_o_sign_lpi_1_dfm_3_mx0c2 = or_181_cse & and_dcpl_1208;
  assign nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_4_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_5_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_6_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_o_mant_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6})
      + conv_u2u_10_11(~ FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6) + 11'b1;
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_7_is_a_greater_oif_aelse_acc_3_nl));
  assign m_row3_4_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10 = ~(m_row2_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row3_3_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10 = ~(m_row2_3_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row3_2_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10 = ~(m_row2_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row3_1_FpAdd_6U_10U_3_a_int_mant_p1_conc_2_10 = ~(m_row2_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row2_4_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10 = ~(m_row1_4_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row2_3_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10 = ~(m_row1_3_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row2_2_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10 = ~(m_row1_2_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign m_row2_1_FpAdd_6U_10U_2_a_int_mant_p1_conc_2_10 = ~(m_row1_1_IsZero_6U_10U_3_aif_IsZero_6U_10U_3_aelse_nor_2
      & (~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000))));
  assign chn_data_in_rsci_oswt_unreg = or_tmp_1099;
  assign chn_data_out_rsci_oswt_unreg = chn_data_out_rsci_bawt & reg_chn_data_out_rsci_ld_core_psct_cse;
  assign IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse = (fsm_output[1]) & (cfg_precision[0]);
  assign FpAdd_6U_10U_7_if_2_and_tmp = (fsm_output[1]) & o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4;
  assign FpAdd_6U_10U_7_if_2_and_tmp_1 = (fsm_output[1]) & reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_7_if_2_and_tmp_2 = (fsm_output[1]) & reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_7_if_2_and_tmp_3 = (fsm_output[1]) & reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_6_if_2_and_tmp = (fsm_output[1]) & reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_6_if_2_and_tmp_1 = (fsm_output[1]) & reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_6_if_2_and_tmp_2 = (fsm_output[1]) & reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_6_if_2_and_tmp_3 = (fsm_output[1]) & o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4;
  assign FpAdd_6U_10U_5_if_2_and_tmp = (fsm_output[1]) & o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  assign FpAdd_6U_10U_5_if_2_and_tmp_1 = (fsm_output[1]) & reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse;
  assign FpAdd_6U_10U_5_if_2_and_tmp_2 = (fsm_output[1]) & o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  assign FpAdd_6U_10U_5_if_2_and_tmp_3 = (fsm_output[1]) & o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4;
  assign FpAdd_6U_10U_4_if_2_and_tmp = (fsm_output[1]) & reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_4_if_2_and_tmp_1 = (fsm_output[1]) & reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_4_if_2_and_tmp_2 = (fsm_output[1]) & reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  assign FpAdd_6U_10U_4_if_2_and_tmp_3 = (fsm_output[1]) & reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_in_rsci_iswt0 <= 1'b0;
      chn_data_out_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_data_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_data_out_rsci_iswt0 <= and_dcpl_66;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_data_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_data_in_rsci_ld_core_psct <= chn_data_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_data_out_rsci_d_0 <= 1'b0;
      chn_data_out_rsci_d_6_1 <= 6'b0;
      chn_data_out_rsci_d_9_7 <= 3'b0;
      chn_data_out_rsci_d_13_10 <= 4'b0;
      chn_data_out_rsci_d_14 <= 1'b0;
      chn_data_out_rsci_d_15 <= 1'b0;
      chn_data_out_rsci_d_16 <= 1'b0;
      chn_data_out_rsci_d_22_17 <= 6'b0;
      chn_data_out_rsci_d_25_23 <= 3'b0;
      chn_data_out_rsci_d_29_26 <= 4'b0;
      chn_data_out_rsci_d_30 <= 1'b0;
      chn_data_out_rsci_d_31 <= 1'b0;
      chn_data_out_rsci_d_32 <= 1'b0;
      chn_data_out_rsci_d_38_33 <= 6'b0;
      chn_data_out_rsci_d_41_39 <= 3'b0;
      chn_data_out_rsci_d_45_42 <= 4'b0;
      chn_data_out_rsci_d_46 <= 1'b0;
      chn_data_out_rsci_d_47 <= 1'b0;
      chn_data_out_rsci_d_48 <= 1'b0;
      chn_data_out_rsci_d_54_49 <= 6'b0;
      chn_data_out_rsci_d_57_55 <= 3'b0;
      chn_data_out_rsci_d_61_58 <= 4'b0;
      chn_data_out_rsci_d_62 <= 1'b0;
      chn_data_out_rsci_d_63 <= 1'b0;
      chn_data_out_rsci_d_64 <= 1'b0;
      chn_data_out_rsci_d_70_65 <= 6'b0;
      chn_data_out_rsci_d_73_71 <= 3'b0;
      chn_data_out_rsci_d_77_74 <= 4'b0;
      chn_data_out_rsci_d_78 <= 1'b0;
      chn_data_out_rsci_d_79 <= 1'b0;
      chn_data_out_rsci_d_80 <= 1'b0;
      chn_data_out_rsci_d_86_81 <= 6'b0;
      chn_data_out_rsci_d_89_87 <= 3'b0;
      chn_data_out_rsci_d_93_90 <= 4'b0;
      chn_data_out_rsci_d_94 <= 1'b0;
      chn_data_out_rsci_d_95 <= 1'b0;
      chn_data_out_rsci_d_96 <= 1'b0;
      chn_data_out_rsci_d_102_97 <= 6'b0;
      chn_data_out_rsci_d_105_103 <= 3'b0;
      chn_data_out_rsci_d_109_106 <= 4'b0;
      chn_data_out_rsci_d_110 <= 1'b0;
      chn_data_out_rsci_d_111 <= 1'b0;
      chn_data_out_rsci_d_112 <= 1'b0;
      chn_data_out_rsci_d_118_113 <= 6'b0;
      chn_data_out_rsci_d_121_119 <= 3'b0;
      chn_data_out_rsci_d_125_122 <= 4'b0;
      chn_data_out_rsci_d_126 <= 1'b0;
      chn_data_out_rsci_d_127 <= 1'b0;
      chn_data_out_rsci_d_128 <= 1'b0;
      chn_data_out_rsci_d_134_129 <= 6'b0;
      chn_data_out_rsci_d_137_135 <= 3'b0;
      chn_data_out_rsci_d_141_138 <= 4'b0;
      chn_data_out_rsci_d_142 <= 1'b0;
      chn_data_out_rsci_d_143 <= 1'b0;
      chn_data_out_rsci_d_144 <= 1'b0;
      chn_data_out_rsci_d_150_145 <= 6'b0;
      chn_data_out_rsci_d_153_151 <= 3'b0;
      chn_data_out_rsci_d_157_154 <= 4'b0;
      chn_data_out_rsci_d_158 <= 1'b0;
      chn_data_out_rsci_d_159 <= 1'b0;
      chn_data_out_rsci_d_160 <= 1'b0;
      chn_data_out_rsci_d_166_161 <= 6'b0;
      chn_data_out_rsci_d_169_167 <= 3'b0;
      chn_data_out_rsci_d_173_170 <= 4'b0;
      chn_data_out_rsci_d_174 <= 1'b0;
      chn_data_out_rsci_d_175 <= 1'b0;
      chn_data_out_rsci_d_176 <= 1'b0;
      chn_data_out_rsci_d_182_177 <= 6'b0;
      chn_data_out_rsci_d_185_183 <= 3'b0;
      chn_data_out_rsci_d_189_186 <= 4'b0;
      chn_data_out_rsci_d_190 <= 1'b0;
      chn_data_out_rsci_d_191 <= 1'b0;
      chn_data_out_rsci_d_192 <= 1'b0;
      chn_data_out_rsci_d_198_193 <= 6'b0;
      chn_data_out_rsci_d_201_199 <= 3'b0;
      chn_data_out_rsci_d_205_202 <= 4'b0;
      chn_data_out_rsci_d_206 <= 1'b0;
      chn_data_out_rsci_d_207 <= 1'b0;
      chn_data_out_rsci_d_208 <= 1'b0;
      chn_data_out_rsci_d_214_209 <= 6'b0;
      chn_data_out_rsci_d_217_215 <= 3'b0;
      chn_data_out_rsci_d_221_218 <= 4'b0;
      chn_data_out_rsci_d_222 <= 1'b0;
      chn_data_out_rsci_d_223 <= 1'b0;
      chn_data_out_rsci_d_224 <= 1'b0;
      chn_data_out_rsci_d_230_225 <= 6'b0;
      chn_data_out_rsci_d_233_231 <= 3'b0;
      chn_data_out_rsci_d_237_234 <= 4'b0;
      chn_data_out_rsci_d_238 <= 1'b0;
      chn_data_out_rsci_d_239 <= 1'b0;
      chn_data_out_rsci_d_240 <= 1'b0;
      chn_data_out_rsci_d_246_241 <= 6'b0;
      chn_data_out_rsci_d_249_247 <= 3'b0;
      chn_data_out_rsci_d_253_250 <= 4'b0;
      chn_data_out_rsci_d_254 <= 1'b0;
      chn_data_out_rsci_d_255 <= 1'b0;
    end
    else if ( chn_data_out_and_cse ) begin
      chn_data_out_rsci_d_0 <= MUX1HOT_s_1_3_2(data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_6_1 <= MUX1HOT_v_6_3_2(o_data_data_0_6_1_sva_10, o_data_data_0_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_9_7 <= MUX1HOT_v_3_3_2(o_data_data_0_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_13_10 <= MUX1HOT_v_4_3_2(o_data_data_0_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_1_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_14 <= MUX1HOT_s_1_3_2(data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_15 <= data_truncate_mux1h_320_itm_4;
      chn_data_out_rsci_d_16 <= MUX1HOT_s_1_3_2(data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_22_17 <= MUX1HOT_v_6_3_2(o_data_data_1_6_1_sva_10, o_data_data_1_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_25_23 <= MUX1HOT_v_3_3_2(o_data_data_1_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_29_26 <= MUX1HOT_v_4_3_2(o_data_data_1_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_3_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_30 <= MUX1HOT_s_1_3_2(data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_2_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_31 <= data_truncate_mux1h_326_itm_4;
      chn_data_out_rsci_d_32 <= MUX1HOT_s_1_3_2(data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_38_33 <= MUX1HOT_v_6_3_2(o_data_data_2_6_1_sva_10, o_data_data_2_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_41_39 <= MUX1HOT_v_3_3_2(o_data_data_2_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_45_42 <= MUX1HOT_v_4_3_2(o_data_data_2_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_5_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_46 <= MUX1HOT_s_1_3_2(data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_4_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_47 <= data_truncate_mux1h_332_itm_4;
      chn_data_out_rsci_d_48 <= MUX1HOT_s_1_3_2(data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_54_49 <= MUX1HOT_v_6_3_2(o_data_data_3_6_1_sva_10, o_data_data_3_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_57_55 <= MUX1HOT_v_3_3_2(o_data_data_3_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_61_58 <= MUX1HOT_v_4_3_2(o_data_data_3_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_7_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_62 <= MUX1HOT_s_1_3_2(data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_6_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_63 <= data_truncate_mux1h_338_itm_4;
      chn_data_out_rsci_d_64 <= MUX1HOT_s_1_3_2(data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_70_65 <= MUX1HOT_v_6_3_2(o_data_data_4_6_1_sva_10, o_data_data_4_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_73_71 <= MUX1HOT_v_3_3_2(o_data_data_4_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_77_74 <= MUX1HOT_v_4_3_2(o_data_data_4_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_9_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_78 <= MUX1HOT_s_1_3_2(data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_8_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_79 <= data_truncate_mux1h_344_itm_4;
      chn_data_out_rsci_d_80 <= MUX1HOT_s_1_3_2(data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_86_81 <= MUX1HOT_v_6_3_2(o_data_data_5_6_1_sva_10, o_data_data_5_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_89_87 <= MUX1HOT_v_3_3_2(o_data_data_5_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_93_90 <= MUX1HOT_v_4_3_2(o_data_data_5_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_11_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_94 <= MUX1HOT_s_1_3_2(data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_10_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_95 <= data_truncate_mux1h_350_itm_4;
      chn_data_out_rsci_d_96 <= MUX1HOT_s_1_3_2(data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_102_97 <= MUX1HOT_v_6_3_2(o_data_data_6_6_1_sva_10, o_data_data_6_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_105_103 <= MUX1HOT_v_3_3_2(o_data_data_6_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_109_106 <= MUX1HOT_v_4_3_2(o_data_data_6_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_13_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_110 <= MUX1HOT_s_1_3_2(data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_12_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_111 <= data_truncate_mux1h_356_itm_4;
      chn_data_out_rsci_d_112 <= MUX1HOT_s_1_3_2(data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_118_113 <= MUX1HOT_v_6_3_2(o_data_data_7_6_1_sva_10, o_data_data_7_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_121_119 <= MUX1HOT_v_3_3_2(o_data_data_7_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_125_122 <= MUX1HOT_v_4_3_2(o_data_data_7_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_15_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_126 <= MUX1HOT_s_1_3_2(data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_14_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_127 <= data_truncate_mux1h_362_itm_4;
      chn_data_out_rsci_d_128 <= MUX1HOT_s_1_3_2(data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_134_129 <= MUX1HOT_v_6_3_2(o_data_data_8_6_1_sva_10, o_data_data_8_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_137_135 <= MUX1HOT_v_3_3_2(o_data_data_8_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_141_138 <= MUX1HOT_v_4_3_2(o_data_data_8_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_17_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_142 <= MUX1HOT_s_1_3_2(data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_16_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_143 <= data_truncate_mux1h_368_itm_4;
      chn_data_out_rsci_d_144 <= MUX1HOT_s_1_3_2(data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_150_145 <= MUX1HOT_v_6_3_2(o_data_data_9_6_1_sva_10, o_data_data_9_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_153_151 <= MUX1HOT_v_3_3_2(o_data_data_9_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_157_154 <= MUX1HOT_v_4_3_2(o_data_data_9_13_10_sva_6, ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_19_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_158 <= MUX1HOT_s_1_3_2(data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_18_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_159 <= data_truncate_mux1h_374_itm_4;
      chn_data_out_rsci_d_160 <= MUX1HOT_s_1_3_2(data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_166_161 <= MUX1HOT_v_6_3_2(o_data_data_10_6_1_sva_10, o_data_data_10_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_169_167 <= MUX1HOT_v_3_3_2(o_data_data_10_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_173_170 <= MUX1HOT_v_4_3_2(o_data_data_10_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_21_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_174 <= MUX1HOT_s_1_3_2(data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_20_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_175 <= data_truncate_mux1h_380_itm_4;
      chn_data_out_rsci_d_176 <= MUX1HOT_s_1_3_2(data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_182_177 <= MUX1HOT_v_6_3_2(o_data_data_11_6_1_sva_10, o_data_data_11_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_185_183 <= MUX1HOT_v_3_3_2(o_data_data_11_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_189_186 <= MUX1HOT_v_4_3_2(o_data_data_11_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_23_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_190 <= MUX1HOT_s_1_3_2(data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_22_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_191 <= data_truncate_mux1h_386_itm_4;
      chn_data_out_rsci_d_192 <= MUX1HOT_s_1_3_2(data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_198_193 <= MUX1HOT_v_6_3_2(o_data_data_12_6_1_sva_10, o_data_data_12_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_201_199 <= MUX1HOT_v_3_3_2(o_data_data_12_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_205_202 <= MUX1HOT_v_4_3_2(o_data_data_12_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_25_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_206 <= MUX1HOT_s_1_3_2(data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_24_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_207 <= data_truncate_mux1h_392_itm_4;
      chn_data_out_rsci_d_208 <= MUX1HOT_s_1_3_2(data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_214_209 <= MUX1HOT_v_6_3_2(o_data_data_13_6_1_sva_10, o_data_data_13_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_217_215 <= MUX1HOT_v_3_3_2(o_data_data_13_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_221_218 <= MUX1HOT_v_4_3_2(o_data_data_13_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_27_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_222 <= MUX1HOT_s_1_3_2(data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_26_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_223 <= data_truncate_mux1h_398_itm_4;
      chn_data_out_rsci_d_224 <= MUX1HOT_s_1_3_2(data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_230_225 <= MUX1HOT_v_6_3_2(o_data_data_14_6_1_sva_10, o_data_data_14_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_233_231 <= MUX1HOT_v_3_3_2(o_data_data_14_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_237_234 <= MUX1HOT_v_4_3_2(o_data_data_14_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_29_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_238 <= MUX1HOT_s_1_3_2(data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_28_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_239 <= data_truncate_mux1h_404_itm_4;
      chn_data_out_rsci_d_240 <= MUX1HOT_s_1_3_2(data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4,
          data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0[0]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_246_241 <= MUX1HOT_v_6_3_2(o_data_data_15_6_1_sva_10, o_data_data_15_6_1_sva_8,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0[6:1]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_249_247 <= MUX1HOT_v_3_3_2(o_data_data_15_9_7_sva_6, ({{2{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0[9:7]), {data_truncate_nor_dfs_4
          , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_253_250 <= MUX1HOT_v_4_3_2(o_data_data_15_13_10_sva_6,
          ({{3{IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}},
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4}),
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_31_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_254 <= MUX1HOT_s_1_3_2(data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4,
          IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4,
          (FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_30_nl),
          {data_truncate_nor_dfs_4 , data_truncate_equal_tmp_4 , data_truncate_nor_tmp_5});
      chn_data_out_rsci_d_255 <= data_truncate_mux1h_410_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_data_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_66 | and_dcpl_68) ) begin
      reg_chn_data_out_rsci_ld_core_psct_cse <= ~ and_dcpl_68;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_1099 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_358_rgt | and_360_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm,
          {and_358_rgt , and_360_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_370_rgt | and_374_rgt | and_dcpl_78 | and_383_rgt |
        and_386_rgt) & (mux_54_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[137:128]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[9:0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w4,
          {and_370_rgt , and_374_rgt , and_dcpl_78 , and_383_rgt , and_386_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_104 | and_388_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp,
          IsNaN_6U_10U_1_land_1_lpi_1_dfm, and_388_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_390_rgt | and_392_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm,
          {and_390_rgt , and_392_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_401_rgt | and_404_rgt | and_dcpl_78 | and_413_rgt |
        and_416_rgt) & (mux_59_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[153:144]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[25:16]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_2_mx0w4,
          {and_401_rgt , and_404_rgt , and_dcpl_78 , and_413_rgt , and_416_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_134 | and_418_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp,
          IsNaN_6U_10U_1_land_2_lpi_1_dfm, and_418_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_420_rgt | and_422_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm,
          {and_420_rgt , and_422_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_431_rgt | and_434_rgt | and_dcpl_78 | and_443_rgt |
        and_446_rgt) & (mux_64_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[169:160]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[41:32]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w4,
          {and_431_rgt , and_434_rgt , and_dcpl_78 , and_443_rgt , and_446_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_164 | and_448_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp,
          IsNaN_6U_10U_1_land_3_lpi_1_dfm, and_448_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_450_rgt | and_452_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_qr_3_0_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_lpi_1_dfm,
          {and_450_rgt , and_452_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_454_rgt | and_456_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm,
          {and_454_rgt , and_456_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_175 | and_459_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp,
          IsNaN_6U_10U_3_land_1_lpi_1_dfm, and_459_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_461_rgt | and_463_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm,
          {and_461_rgt , and_463_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_182 | and_466_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp,
          IsNaN_6U_10U_3_land_2_lpi_1_dfm, and_466_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_468_rgt | and_470_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm,
          {and_468_rgt , and_470_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_189 | and_473_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp,
          IsNaN_6U_10U_3_land_3_lpi_1_dfm, and_473_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_475_rgt | and_477_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm,
          {and_475_rgt , and_477_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_479_rgt | and_481_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm,
          {and_479_rgt , and_481_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_200 | and_484_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp,
          IsNaN_6U_10U_5_land_1_lpi_1_dfm, and_484_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_486_rgt | and_488_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm,
          {and_486_rgt , and_488_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_207 | and_491_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp,
          IsNaN_6U_10U_5_land_2_lpi_1_dfm, and_491_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_493_rgt | and_495_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm,
          {and_493_rgt , and_495_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_214 | and_498_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp,
          IsNaN_6U_10U_5_land_3_lpi_1_dfm, and_498_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_500_rgt | and_502_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm,
          {and_500_rgt , and_502_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_504_rgt | and_506_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm,
          {and_504_rgt , and_506_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_225 | and_509_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp,
          IsNaN_6U_10U_7_land_1_lpi_1_dfm, and_509_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_511_rgt | and_513_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm,
          {and_511_rgt , and_513_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_232 | and_516_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp,
          IsNaN_6U_10U_7_land_2_lpi_1_dfm, and_516_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_518_rgt | and_520_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm,
          {and_518_rgt , and_520_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_239 | and_523_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp,
          IsNaN_6U_10U_7_land_3_lpi_1_dfm, and_523_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( core_wen & (and_525_rgt | and_527_rgt | and_dcpl_78) & mux_tmp_49 )
        begin
      FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_3 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm,
          {and_525_rgt , and_527_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse <= 1'b0;
      reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_4_land_lpi_1_dfm_st_2 <= 1'b0;
      reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_4_land_3_lpi_1_dfm_3 <= 1'b0;
      reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_4_land_2_lpi_1_dfm_3 <= 1'b0;
      reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_4_land_1_lpi_1_dfm_3 <= 1'b0;
      reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_2 <= 1'b0;
      reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_3 <= 1'b0;
      reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_3 <= 1'b0;
      reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_3 <= 1'b0;
      reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse <= 1'b0;
      reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= 1'b0;
      reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse <= 1'b0;
      reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= 1'b0;
      o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= 1'b0;
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= 1'b0;
      o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= 1'b0;
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= 1'b0;
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= 1'b0;
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= 1'b0;
      IntSubExt_16U_16U_17U_2_o_acc_2_itm_2 <= 17'b0;
      m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2 <= 17'b0;
      IntSubExt_16U_16U_17U_1_o_acc_2_itm_2 <= 17'b0;
      m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2 <= 17'b0;
      IntAddExt_16U_16U_17U_o_acc_1_itm_2 <= 17'b0;
      m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2 <= 17'b0;
      IntSubExt_16U_16U_17U_o_acc_2_itm_2 <= 17'b0;
      m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2 <= 17'b0;
      m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2 <= 17'b0;
      m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2 <= 17'b0;
      m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2 <= 17'b0;
      m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2 <= 17'b0;
      IntSubExt_16U_16U_17U_2_o_acc_1_itm_2 <= 17'b0;
      IntSubExt_16U_16U_17U_1_o_acc_1_itm_2 <= 17'b0;
      IntAddExt_16U_16U_17U_o_acc_itm_2 <= 17'b0;
      IntSubExt_16U_16U_17U_o_acc_1_itm_2 <= 17'b0;
    end
    else if ( IsNaN_6U_10U_6_aelse_and_8_cse ) begin
      reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp,
          IsNaN_6U_10U_6_land_lpi_1_dfm_st, and_dcpl_78);
      reg_m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0,
          m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp,
          IsNaN_6U_10U_6_land_3_lpi_1_dfm, and_dcpl_78);
      reg_m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0,
          m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp,
          IsNaN_6U_10U_6_land_2_lpi_1_dfm, and_dcpl_78);
      reg_m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0,
          m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp,
          IsNaN_6U_10U_6_land_1_lpi_1_dfm, and_dcpl_78);
      reg_m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0,
          m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_4_land_lpi_1_dfm_st_2 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp,
          IsNaN_6U_10U_4_land_lpi_1_dfm_st, and_dcpl_78);
      reg_m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0,
          m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_4_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp,
          IsNaN_6U_10U_4_land_3_lpi_1_dfm, and_dcpl_78);
      reg_m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0,
          m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_4_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp,
          IsNaN_6U_10U_4_land_2_lpi_1_dfm, and_dcpl_78);
      reg_m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0,
          m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_4_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp,
          IsNaN_6U_10U_4_land_1_lpi_1_dfm, and_dcpl_78);
      reg_m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0,
          m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_2 <= MUX_s_1_2_2(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp,
          IsNaN_6U_10U_2_land_lpi_1_dfm_st, and_dcpl_78);
      reg_m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= MUX_s_1_2_2(m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp,
          IsNaN_6U_10U_2_land_3_lpi_1_dfm, and_dcpl_78);
      reg_m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= MUX_s_1_2_2(m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp,
          IsNaN_6U_10U_2_land_2_lpi_1_dfm, and_dcpl_78);
      reg_m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= MUX_s_1_2_2(m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st,
          and_dcpl_78);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp,
          IsNaN_6U_10U_2_land_1_lpi_1_dfm, and_dcpl_78);
      reg_m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_1_cse
          <= MUX_s_1_2_2(m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp,
          IsNaN_6U_10U_land_lpi_1_dfm_st, and_dcpl_78);
      reg_m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0,
          m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp,
          IsNaN_6U_10U_land_3_lpi_1_dfm, and_dcpl_78);
      reg_m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0,
          m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp,
          IsNaN_6U_10U_land_2_lpi_1_dfm, and_dcpl_78);
      reg_m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0,
          m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st,
          and_dcpl_78);
      reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_and_tmp,
          IsNaN_6U_10U_land_1_lpi_1_dfm, and_dcpl_78);
      reg_m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_1_cse
          <= MUX_s_1_2_2(m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0,
          m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0,
          o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0,
          o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0,
          o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0,
          o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= MUX_s_1_2_2(o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0,
          o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st,
          and_dcpl_78);
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= MUX_s_1_2_2(o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0,
          o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st,
          and_dcpl_78);
      o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= MUX_s_1_2_2(o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0,
          o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st,
          and_dcpl_78);
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3
          <= MUX_s_1_2_2(o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0,
          o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st,
          and_dcpl_78);
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0,
          o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0,
          o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0,
          o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0,
          o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0,
          o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0,
          o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0,
          o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st,
          and_dcpl_78);
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3
          <= MUX_s_1_2_2(o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0,
          o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st,
          and_dcpl_78);
      IntSubExt_16U_16U_17U_2_o_acc_2_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0,
          IntSubExt_16U_16U_17U_2_o_acc_2_itm, and_dcpl_245);
      m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0,
          m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva, and_dcpl_245);
      IntSubExt_16U_16U_17U_1_o_acc_2_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0,
          IntSubExt_16U_16U_17U_1_o_acc_2_itm, and_dcpl_245);
      m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0,
          m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva, and_dcpl_245);
      IntAddExt_16U_16U_17U_o_acc_1_itm_2 <= MUX_v_17_2_2(IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0,
          IntAddExt_16U_16U_17U_o_acc_1_itm, and_dcpl_245);
      m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0,
          m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva, and_dcpl_245);
      IntSubExt_16U_16U_17U_o_acc_2_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0,
          IntSubExt_16U_16U_17U_o_acc_2_itm, and_dcpl_245);
      m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0,
          m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva, and_dcpl_245);
      m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0,
          m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva, and_dcpl_245);
      m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0,
          m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva, and_dcpl_245);
      m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0,
          m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva, and_dcpl_245);
      m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_2 <= MUX_v_17_2_2(m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0,
          m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva, and_dcpl_245);
      IntSubExt_16U_16U_17U_2_o_acc_1_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0,
          IntSubExt_16U_16U_17U_2_o_acc_1_itm, and_dcpl_245);
      IntSubExt_16U_16U_17U_1_o_acc_1_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0,
          IntSubExt_16U_16U_17U_1_o_acc_1_itm, and_dcpl_245);
      IntAddExt_16U_16U_17U_o_acc_itm_2 <= MUX_v_17_2_2(IntAddExt_16U_16U_17U_o_acc_itm_mx0w0,
          IntAddExt_16U_16U_17U_o_acc_itm, and_dcpl_245);
      IntSubExt_16U_16U_17U_o_acc_1_itm_2 <= MUX_v_17_2_2(IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0,
          IntSubExt_16U_16U_17U_o_acc_1_itm, and_dcpl_245);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_a_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_a_int_mant_p1_and_cse ) begin
      FpAdd_6U_10U_3_a_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_3_a_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_3_b_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_3_b_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp,
          FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_1, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_537_rgt | and_540_rgt | and_dcpl_78 | and_548_rgt |
        and_551_rgt) & (mux_72_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[105:96]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[233:224]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_4_mx0w4,
          {and_537_rgt , and_540_rgt , and_dcpl_78 , and_548_rgt , and_551_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_3_mx0[1]),
          {and_dcpl_269 , and_dcpl_270 , and_dcpl_271});
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_0_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_3_mx0[0]),
          {and_dcpl_269 , and_dcpl_270 , and_dcpl_271});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_269 | and_dcpl_78 | and_dcpl_239) & mux_tmp_76
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2,
          {and_dcpl_269 , and_dcpl_78 , and_dcpl_239});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_a_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_a_int_mant_p1_and_7_cse ) begin
      FpAdd_6U_10U_3_a_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_3_a_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_3_b_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_3_b_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp,
          FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_3_a_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_3_a_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_3_b_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_3_b_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp,
          FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_3_a_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_a_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_3_a_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_3_b_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_3_b_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_3_b_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp,
          FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_2_a_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_2_a_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_2_b_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_2_b_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp,
          FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_2_a_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_2_a_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_2_b_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_2_b_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp,
          FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_2_a_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_2_a_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_2_b_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_2_b_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp,
          FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_2_a_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_a_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_2_a_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_2_b_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_2_b_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_2_b_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp,
          FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_1_a_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_1_a_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_1_b_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp,
          FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_1_a_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_1_a_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_1_b_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp,
          FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_1_a_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_1_a_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_1_b_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp,
          FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_a_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_a_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_b_int_mant_p1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_sva_mx0w0,
          FpAdd_6U_10U_b_int_mant_p1_sva, and_dcpl_78);
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp,
          FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_a_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_3_sva_mx0w0,
          FpAdd_6U_10U_b_int_mant_p1_3_sva, and_dcpl_78);
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp,
          FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_a_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_b_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp,
          FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1, and_dcpl_78);
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_a_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_1_sva_mx0w0,
          FpAdd_6U_10U_b_int_mant_p1_1_sva, and_dcpl_78);
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp,
          FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_564_rgt | and_567_rgt | and_dcpl_78 | and_575_rgt |
        and_578_rgt) & (mux_84_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[89:80]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[217:208]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_2_mx0w4,
          {and_564_rgt , and_567_rgt , and_dcpl_78 , and_575_rgt , and_578_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_3_mx0[1]),
          {and_dcpl_295 , and_dcpl_296 , and_dcpl_297});
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_0_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_3_mx0[0]),
          {and_dcpl_295 , and_dcpl_296 , and_dcpl_297});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_295 | and_dcpl_78 | and_dcpl_232) & mux_tmp_88
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2,
          {and_dcpl_295 , and_dcpl_78 , and_dcpl_232});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_590_rgt | and_593_rgt | and_dcpl_78 | and_601_rgt |
        and_604_rgt) & (mux_96_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[73:64]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[201:192]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_mx0w4,
          {and_590_rgt , and_593_rgt , and_dcpl_78 , and_601_rgt , and_604_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_3_mx0[1]),
          {and_dcpl_321 , and_dcpl_322 , and_dcpl_323});
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_0_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_3_mx0[0]),
          {and_dcpl_321 , and_dcpl_322 , and_dcpl_323});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_321 | and_dcpl_78 | and_dcpl_225) & mux_tmp_100
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2,
          {and_dcpl_321 , and_dcpl_78 , and_dcpl_225});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_610_rgt | and_612_rgt | and_dcpl_78 | and_614_rgt |
        and_616_rgt) & (mux_108_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[169:160]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[105:96]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          {and_610_rgt , and_612_rgt , and_dcpl_78 , and_614_rgt , and_616_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_7 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          {and_dcpl_333 , and_dcpl_78 , and_dcpl_214});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          {and_dcpl_333 , and_dcpl_78 , and_dcpl_214});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          {and_dcpl_333 , and_dcpl_78 , and_dcpl_214});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_620_rgt | and_622_rgt | and_dcpl_78 | and_624_rgt |
        and_626_rgt) & (mux_117_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[153:144]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[89:80]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          {and_620_rgt , and_622_rgt , and_dcpl_78 , and_624_rgt , and_626_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_7 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          {and_dcpl_343 , and_dcpl_78 , and_dcpl_207});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          {and_dcpl_343 , and_dcpl_78 , and_dcpl_207});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          {and_dcpl_343 , and_dcpl_78 , and_dcpl_207});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_630_rgt | and_632_rgt | and_dcpl_78 | and_634_rgt |
        and_636_rgt) & (mux_126_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[137:128]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[73:64]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          {and_630_rgt , and_632_rgt , and_dcpl_78 , and_634_rgt , and_636_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_7 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          {and_dcpl_353 , and_dcpl_78 , and_dcpl_200});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          {and_dcpl_353 , and_dcpl_78 , and_dcpl_200});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          {and_dcpl_353 , and_dcpl_78 , and_dcpl_200});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_640_rgt | and_642_rgt | and_dcpl_78 | and_644_rgt |
        and_646_rgt) & (mux_138_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[105:96]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[169:160]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          {and_640_rgt , and_642_rgt , and_dcpl_78 , and_644_rgt , and_646_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]), FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1_1,
          {and_dcpl_363 , and_dcpl_189 , and_dcpl_364});
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_mx0[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_1, {and_dcpl_363
          , and_dcpl_189 , and_dcpl_364});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_649_rgt | and_dcpl_78 | and_dcpl_189) & mux_tmp_142
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          {and_649_rgt , and_dcpl_78 , and_dcpl_189});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_652_rgt | and_654_rgt | and_dcpl_78 | and_656_rgt |
        and_658_rgt) & (mux_147_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[89:80]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[153:144]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          {and_652_rgt , and_654_rgt , and_dcpl_78 , and_656_rgt , and_658_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]), FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1_1,
          {and_dcpl_375 , and_dcpl_182 , and_dcpl_376});
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_mx0[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_1, {and_dcpl_375
          , and_dcpl_182 , and_dcpl_376});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_661_rgt | and_dcpl_78 | and_dcpl_182) & mux_tmp_151
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          {and_661_rgt , and_dcpl_78 , and_dcpl_182});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_a_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_a_int_mant_p1_and_8_cse ) begin
      FpAdd_6U_10U_1_a_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_a_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_1_a_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2 <= MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_2_sva_mx0w0,
          FpAdd_6U_10U_1_b_int_mant_p1_2_sva, and_dcpl_78);
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_4 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp,
          FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_664_rgt | and_666_rgt | and_dcpl_78 | and_668_rgt |
        and_670_rgt) & (mux_158_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[73:64]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[137:128]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          {and_664_rgt , and_666_rgt , and_dcpl_78 , and_668_rgt , and_670_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]), FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1_1,
          {and_dcpl_387 , and_dcpl_175 , and_dcpl_388});
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_mx0[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_1, {and_dcpl_387
          , and_dcpl_175 , and_dcpl_388});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_673_rgt | and_dcpl_78 | and_dcpl_175) & mux_tmp_162
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          {and_673_rgt , and_dcpl_78 , and_dcpl_175});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_mx0[1]), and_dcpl_391);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5_0_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_mx0[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_mx0[0]), and_dcpl_391);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_164 | and_dcpl_78 | and_676_rgt) & mux_tmp_172
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2,
          {and_dcpl_164 , and_dcpl_78 , and_676_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_mx0[1]), and_dcpl_394);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5_0_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_mx0[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_mx0[0]), and_dcpl_394);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_134 | and_dcpl_78 | and_680_rgt) & mux_tmp_179
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2,
          {and_dcpl_134 , and_dcpl_78 , and_680_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_mx0[1]), and_dcpl_397);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5_0_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_mx0[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_mx0[0]), and_dcpl_397);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_104 | and_dcpl_78 | and_683_rgt) & mux_tmp_186
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2,
          {and_dcpl_104 , and_dcpl_78 , and_683_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_tmp_56 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_land_1_lpi_1_dfm_2_cse)
        | and_689_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_7,
          FpAdd_6U_10U_FpAdd_6U_10U_or_4_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_13_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_land_3_lpi_1_dfm_2_cse)
        | and_691_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_7,
          FpAdd_6U_10U_FpAdd_6U_10U_or_6_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_12_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_2_land_1_lpi_1_dfm_3) | and_693_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_7,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_4_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_13_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_2_land_3_lpi_1_dfm_3) | and_695_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_6_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_12_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_land_1_lpi_1_dfm_3) | and_697_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_7,
          FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_4_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_13_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_land_3_lpi_1_dfm_3) | and_699_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_7,
          FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_6_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_12_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_6_land_1_lpi_1_dfm_2_cse)
        | and_701_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_7,
          FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_4_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_13_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_6_land_3_lpi_1_dfm_2_cse)
        | and_703_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_7,
          FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_6_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_12_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_land_2_lpi_1_dfm_2_cse)
        | and_705_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_7,
          FpAdd_6U_10U_FpAdd_6U_10U_or_5_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_11_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_2_land_2_lpi_1_dfm_3) | and_707_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_7,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_5_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_11_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_land_2_lpi_1_dfm_3) | and_709_rgt)
        & mux_468_cse ) begin
      FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_7,
          FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_5_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_11_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((or_181_cse & reg_IsNaN_6U_10U_6_land_2_lpi_1_dfm_2_cse)
        | and_711_rgt) & mux_468_cse ) begin
      FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_7,
          FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_5_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_11_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_713_rgt | and_715_rgt | and_dcpl_78) & mux_468_cse
        ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_FpAdd_6U_10U_or_11_itm, FpAdd_6U_10U_o_mant_lpi_1_dfm_2, {(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_nl)
          , (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_10_nl) , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_717_rgt | and_719_rgt | and_dcpl_78) & mux_468_cse
        ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_11_itm, FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2,
          {(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_nl) , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_10_nl)
          , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_721_rgt | and_723_rgt | and_dcpl_78) & mux_468_cse
        ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_11_itm, FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2,
          {(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_nl) , (FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_10_nl)
          , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_725_rgt | and_727_rgt | and_dcpl_78) & mux_468_cse
        ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_11_itm, FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2,
          {(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_nl) , (FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_10_nl)
          , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4
          <= 1'b0;
      reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4
          <= 1'b0;
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= 1'b0;
      reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse
          <= 1'b0;
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= 1'b0;
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= 1'b0;
      reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= 1'b0;
      IsNaN_6U_10U_15_land_3_lpi_1_dfm_4 <= 1'b0;
      m_row0_unequal_tmp_3 <= 1'b0;
      IsNaN_6U_10U_15_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_15_land_1_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_15_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_12_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_10_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_4 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2 <= 4'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_o_expo_and_cse ) begin
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4
          <= o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
      reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
      reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
      reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse
          <= o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_3;
      reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
      reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
      reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse
          <= o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4
          <= o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_3;
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
      reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse
          <= o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4
          <= o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_3;
      reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
      reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
      reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
      reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse
          <= o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_3;
      IsNaN_6U_10U_15_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_2_tmp;
      m_row0_unequal_tmp_3 <= ~((cfg_precision==2'b10));
      IsNaN_6U_10U_15_land_2_lpi_1_dfm_4 <= IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_1_tmp;
      IsNaN_6U_10U_15_land_1_lpi_1_dfm_4 <= IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_tmp;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp;
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_4 <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_4 <= IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp;
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp;
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp;
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp;
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp;
      IsNaN_6U_10U_15_land_lpi_1_dfm_4 <= IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_3_tmp;
      IsNaN_6U_10U_12_land_lpi_1_dfm_4 <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp;
      IsNaN_6U_10U_10_land_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp;
      IsNaN_6U_10U_8_land_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_3_o_expo_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_2_o_expo_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_o_expo_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp <= FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1 <= FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_4;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2 <= FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_10_land_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_12_land_lpi_1_dfm_st_3 <= 1'b0;
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= 1'b0;
      reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= 1'b0;
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= 1'b0;
      reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= 1'b0;
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= 1'b0;
      reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= 1'b0;
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= 1'b0;
      reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= 1'b0;
      reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse <= 1'b0;
      reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse <= 1'b0;
      reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1 <= 1'b0;
      reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1 <= 1'b0;
      o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= 1'b0;
      o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= 1'b0;
      o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= 1'b0;
      o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_12_aelse_and_4_cse ) begin
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp,
          IsNaN_6U_10U_12_land_2_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp,
          IsNaN_6U_10U_8_land_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp,
          IsNaN_6U_10U_8_land_3_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp,
          IsNaN_6U_10U_8_land_2_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp,
          IsNaN_6U_10U_14_land_1_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp,
          IsNaN_6U_10U_14_land_2_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp,
          IsNaN_6U_10U_14_land_3_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_10_land_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp,
          IsNaN_6U_10U_14_land_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp,
          IsNaN_6U_10U_12_land_1_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp,
          IsNaN_6U_10U_12_land_3_lpi_1_dfm_st, and_dcpl_78);
      IsNaN_6U_10U_12_land_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp,
          IsNaN_6U_10U_12_land_lpi_1_dfm_st, and_dcpl_78);
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= MUX_s_1_2_2(o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0,
          o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm, and_dcpl_78);
      reg_o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= MUX_s_1_2_2(o_col1_4_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0,
          o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm, and_dcpl_78);
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= MUX_s_1_2_2(o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0,
          o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm, and_dcpl_78);
      reg_o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= MUX_s_1_2_2(o_col1_3_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0,
          o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm, and_dcpl_78);
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= MUX_s_1_2_2(o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0,
          o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm, and_dcpl_78);
      reg_o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= MUX_s_1_2_2(o_col1_2_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0,
          o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm, and_dcpl_78);
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_2 <= MUX_s_1_2_2(o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0,
          o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm, and_dcpl_78);
      reg_o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_cse <= MUX_s_1_2_2(o_col1_1_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0,
          o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm, and_dcpl_78);
      reg_o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse <= MUX_s_1_2_2(o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0,
          o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm, and_dcpl_78);
      reg_o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse <= MUX_s_1_2_2(o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0,
          o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm, and_dcpl_78);
      reg_o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1 <= MUX_s_1_2_2(o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0,
          o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm, and_dcpl_78);
      reg_o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_cse_1 <= MUX_s_1_2_2(o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0,
          o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm, and_dcpl_78);
      o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= MUX_s_1_2_2(o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0,
          o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm, and_dcpl_78);
      o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= MUX_s_1_2_2(o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0,
          o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm, and_dcpl_78);
      o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= MUX_s_1_2_2(o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0,
          o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm, and_dcpl_78);
      o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_2 <= MUX_s_1_2_2(o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0,
          o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & main_stage_v_2) | main_stage_v_3_mx0c1) )
        begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_14_land_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_12_land_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 <= 1'b0;
      data_truncate_equal_tmp_3 <= 1'b0;
      data_truncate_nor_tmp_4 <= 1'b0;
      data_truncate_nor_dfs_3 <= 1'b0;
      data_truncate_mux1h_410_itm_3 <= 1'b0;
      data_truncate_mux1h_404_itm_3 <= 1'b0;
      data_truncate_mux1h_398_itm_3 <= 1'b0;
      data_truncate_mux1h_392_itm_3 <= 1'b0;
      data_truncate_mux1h_386_itm_3 <= 1'b0;
      data_truncate_mux1h_380_itm_3 <= 1'b0;
      data_truncate_mux1h_374_itm_3 <= 1'b0;
      data_truncate_mux1h_368_itm_3 <= 1'b0;
      data_truncate_mux1h_362_itm_3 <= 1'b0;
      data_truncate_mux1h_356_itm_3 <= 1'b0;
      data_truncate_mux1h_350_itm_3 <= 1'b0;
      data_truncate_mux1h_344_itm_3 <= 1'b0;
      data_truncate_mux1h_338_itm_3 <= 1'b0;
      data_truncate_mux1h_332_itm_3 <= 1'b0;
      data_truncate_mux1h_326_itm_3 <= 1'b0;
      data_truncate_mux1h_320_itm_3 <= 1'b0;
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_3 <= 1'b0;
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_3 <= 1'b0;
      IsNaN_6U_10U_9_land_lpi_1_dfm_3 <= 1'b0;
      IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_11_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_13_land_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_13_land_2_lpi_1_dfm_3 <= 1'b0;
      IsNaN_6U_10U_13_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_13_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_15_land_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_15_land_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_15_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_15_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_14_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_10_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_5 <= 1'b0;
      m_row0_unequal_tmp_4 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_14_aelse_and_cse ) begin
      IsNaN_6U_10U_14_land_lpi_1_dfm_st_4 <= IsNaN_6U_10U_10_land_lpi_1_dfm_st_3;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_st_4 <= IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_st_4 <= IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_st_4 <= IsNaN_6U_10U_10_land_1_lpi_1_dfm_st_3;
      IsNaN_6U_10U_12_land_lpi_1_dfm_st_4 <= IsNaN_6U_10U_12_land_lpi_1_dfm_st_3;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_4 <= IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_3;
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_4 <= IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_4 <= IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_3;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 <= IsNaN_6U_10U_8_land_lpi_1_dfm_st_3;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 <= IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 <= IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3;
      data_truncate_equal_tmp_3 <= data_truncate_equal_tmp_mx0w0;
      data_truncate_nor_tmp_4 <= data_truncate_nor_tmp_mx0w0;
      data_truncate_nor_dfs_3 <= data_truncate_nor_dfs_mx0w0;
      data_truncate_mux1h_410_itm_3 <= MUX1HOT_s_1_3_2((z_out[17]), FpAdd_6U_10U_7_mux_61_mx1w0,
          FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2, {data_truncate_data_truncate_nor_1_cse
          , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_404_itm_3 <= MUX1HOT_s_1_4_2((z_out_15[17]), (z_out_1[17]),
          FpAdd_6U_10U_6_mux_61_mx1w1, FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_398_itm_3 <= MUX1HOT_s_1_4_2((z_out_14[17]), (z_out_2[17]),
          FpAdd_6U_10U_5_mux_61_mx1w1, FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_392_itm_3 <= MUX1HOT_s_1_4_2((z_out_13[17]), (z_out_3[17]),
          FpAdd_6U_10U_4_mux_61_mx1w1, FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_386_itm_3 <= MUX1HOT_s_1_4_2((z_out_12[17]), (z_out_4[17]),
          FpAdd_6U_10U_7_mux_45_mx1w0, FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_380_itm_3 <= MUX1HOT_s_1_4_2((z_out_11[17]), (z_out_5[17]),
          FpAdd_6U_10U_6_mux_45_mx1w1, FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_374_itm_3 <= MUX1HOT_s_1_4_2((z_out_10[17]), (z_out_6[17]),
          FpAdd_6U_10U_5_mux_45_mx1w1, FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_368_itm_3 <= MUX1HOT_s_1_4_2((z_out_9[17]), (z_out_7[17]),
          FpAdd_6U_10U_4_mux_45_mx1w1, FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_362_itm_3 <= MUX1HOT_s_1_3_2((z_out_8[17]), FpAdd_6U_10U_7_mux_29_mx1w0,
          FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2, {data_truncate_data_truncate_nor_1_cse
          , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_356_itm_3 <= MUX1HOT_s_1_4_2((z_out_7[17]), (z_out_9[17]),
          FpAdd_6U_10U_6_mux_29_mx1w1, FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_350_itm_3 <= MUX1HOT_s_1_4_2((z_out_6[17]), (z_out_10[17]),
          FpAdd_6U_10U_5_mux_29_mx1w1, FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_344_itm_3 <= MUX1HOT_s_1_4_2((z_out_5[17]), (z_out_11[17]),
          FpAdd_6U_10U_4_mux_29_mx1w1, FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_338_itm_3 <= MUX1HOT_s_1_4_2((z_out_4[17]), (z_out_12[17]),
          FpAdd_6U_10U_7_mux_13_mx1w0, FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_332_itm_3 <= MUX1HOT_s_1_4_2((z_out_3[17]), (z_out_13[17]),
          FpAdd_6U_10U_6_mux_13_mx1w1, FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_326_itm_3 <= MUX1HOT_s_1_4_2((z_out_2[17]), (z_out_14[17]),
          FpAdd_6U_10U_5_mux_13_mx1w1, FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      data_truncate_mux1h_320_itm_3 <= MUX1HOT_s_1_4_2((z_out_1[17]), (z_out_15[17]),
          FpAdd_6U_10U_4_mux_13_mx1w1, FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5, {data_truncate_and_124_cse
          , data_truncate_and_125_cse , data_truncate_and_129_cse , data_truncate_and_130_cse});
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_12_land_1_lpi_1_dfm_4;
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_3 <= IsNaN_6U_10U_9_land_2_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_3 <= IsNaN_6U_10U_9_land_3_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_9_land_lpi_1_dfm_3 <= IsNaN_6U_10U_9_land_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 <= IsNaN_6U_10U_12_land_2_lpi_1_dfm_4;
      IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_12_land_3_lpi_1_dfm_4;
      IsNaN_6U_10U_11_land_lpi_1_dfm_5 <= IsNaN_6U_10U_12_land_lpi_1_dfm_4;
      IsNaN_6U_10U_13_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_13_land_1_lpi_1_dfm_4;
      IsNaN_6U_10U_13_land_2_lpi_1_dfm_3 <= nor_384_cse;
      IsNaN_6U_10U_13_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_13_land_3_lpi_1_dfm_4;
      IsNaN_6U_10U_13_land_lpi_1_dfm_5 <= IsNaN_6U_10U_13_land_lpi_1_dfm_4;
      IsNaN_6U_10U_15_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_15_land_1_lpi_1_dfm_4;
      IsNaN_6U_10U_15_land_2_lpi_1_dfm_5 <= IsNaN_6U_10U_15_land_2_lpi_1_dfm_4;
      IsNaN_6U_10U_15_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_15_land_3_lpi_1_dfm_4;
      IsNaN_6U_10U_15_land_lpi_1_dfm_5 <= IsNaN_6U_10U_15_land_lpi_1_dfm_4;
      IsNaN_6U_10U_14_land_lpi_1_dfm_5 <= IsNaN_6U_10U_14_land_lpi_1_dfm_st;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_14_land_3_lpi_1_dfm_st;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_5 <= IsNaN_6U_10U_14_land_2_lpi_1_dfm_st;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_14_land_1_lpi_1_dfm_st;
      IsNaN_6U_10U_10_land_lpi_1_dfm_5 <= IsNaN_6U_10U_10_land_lpi_1_dfm_4;
      IsNaN_6U_10U_10_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_10_land_3_lpi_1_dfm_4;
      IsNaN_6U_10U_10_land_2_lpi_1_dfm_5 <= IsNaN_6U_10U_10_land_2_lpi_1_dfm_4;
      IsNaN_6U_10U_10_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_10_land_1_lpi_1_dfm_4;
      IsNaN_6U_10U_8_land_lpi_1_dfm_5 <= IsNaN_6U_10U_8_land_lpi_1_dfm_4;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_5 <= IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_5 <= IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_5 <= IsNaN_6U_10U_8_land_1_lpi_1_dfm_4;
      m_row0_unequal_tmp_4 <= m_row0_unequal_tmp_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_int_mant_p1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4)))
        & (~(or_181_cse & o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_4))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_7_int_mant_p1_sva_3 <= readslicef_25_24_1((acc_16_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_int_mant_p1_3_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_7_int_mant_p1_3_sva_3 <= readslicef_25_24_1((acc_17_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_int_mant_p1_2_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_7_int_mant_p1_2_sva_3 <= readslicef_25_24_1((acc_18_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_int_mant_p1_1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_7_int_mant_p1_1_sva_3 <= readslicef_25_24_1((acc_19_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_int_mant_p1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_6_int_mant_p1_sva_3 <= readslicef_25_24_1((acc_20_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_int_mant_p1_3_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_6_int_mant_p1_3_sva_3 <= readslicef_25_24_1((acc_21_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_int_mant_p1_2_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_6_int_mant_p1_2_sva_3 <= readslicef_25_24_1((acc_22_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_int_mant_p1_1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4)))
        & (~(or_181_cse & o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st_4))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_6_int_mant_p1_1_sva_3 <= readslicef_25_24_1((acc_23_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_int_mant_p1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4)))
        & (~(or_181_cse & o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_5_int_mant_p1_sva_3 <= readslicef_25_24_1((acc_24_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_int_mant_p1_3_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_5_int_mant_p1_3_sva_3 <= readslicef_25_24_1((acc_25_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_int_mant_p1_2_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4)))
        & (~(or_181_cse & o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_5_int_mant_p1_2_sva_3 <= readslicef_25_24_1((acc_26_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_int_mant_p1_1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4)))
        & (~(or_181_cse & o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st_4))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_5_int_mant_p1_1_sva_3 <= readslicef_25_24_1((acc_27_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_int_mant_p1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_4_int_mant_p1_sva_3 <= readslicef_25_24_1((acc_28_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_int_mant_p1_3_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_4_int_mant_p1_3_sva_3 <= readslicef_25_24_1((acc_29_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_int_mant_p1_2_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_4_int_mant_p1_2_sva_3 <= readslicef_25_24_1((acc_30_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_int_mant_p1_1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_181_cse & (~ reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse)))
        & (~(or_181_cse & reg_o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st_2_cse))))
        & mux_tmp_191 ) begin
      FpAdd_6U_10U_4_int_mant_p1_1_sva_3 <= readslicef_25_24_1((acc_31_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_828_cse | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_200 | data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_200)) ) begin
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_206 | data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_206)) ) begin
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_212 | data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_212)) ) begin
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_218 | data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_218)) ) begin
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_224 | data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_224)) ) begin
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_230 | data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_230)) ) begin
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_236 | data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_236)) ) begin
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_242 | data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_242)) ) begin
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_248 | data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_248)) ) begin
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_254 | data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_254)) ) begin
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_260 | data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_260)) ) begin
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_266 | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_266)) ) begin
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_272 | data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_272)) ) begin
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_278 | data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_278)) ) begin
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_284 | data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_284)) ) begin
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_290 | data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1))
        ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs
          <= data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_290)) ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs
          <= data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_15_lpi_1_dfm_3 <= 1'b0;
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_14_lpi_1_dfm_3 <= 1'b0;
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_12_lpi_1_dfm_3 <= 1'b0;
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_11_lpi_1_dfm_3 <= 1'b0;
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_10_lpi_1_dfm_3 <= 1'b0;
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_9_lpi_1_dfm_3 <= 1'b0;
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_8_lpi_1_dfm_3 <= 1'b0;
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_7_lpi_1_dfm_3 <= 1'b0;
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_6_lpi_1_dfm_3 <= 1'b0;
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_5_lpi_1_dfm_3 <= 1'b0;
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_4_lpi_1_dfm_3 <= 1'b0;
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_3_lpi_1_dfm_3 <= 1'b0;
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_2_lpi_1_dfm_3 <= 1'b0;
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= 1'b0;
      IsNaN_6U_10U_16_land_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_cse ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_15_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_14_tmp;
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_14_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_13_tmp;
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_12_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_11_tmp;
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_11_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_10_tmp;
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_10_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_9_tmp;
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_9_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_8_tmp;
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_8_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_7_tmp;
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_7_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_6_tmp;
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_6_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_5_tmp;
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_5_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_4_tmp;
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_4_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_3_tmp;
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_3_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_2_tmp;
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_2_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_1_tmp;
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
          <= data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_land_1_lpi_1_dfm_3 <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_16_nor_15_itm_2 <= 1'b0;
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm_2 <= 1'b0;
      IsNaN_6U_10U_16_nor_12_itm_2 <= 1'b0;
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_16_and_4_cse ) begin
      IsNaN_6U_10U_16_nor_15_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_16_nor_15_tmp, IsNaN_6U_10U_16_nor_15_itm,
          and_dcpl_547);
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_tmp,
          IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm, and_dcpl_547);
      IsNaN_6U_10U_16_nor_12_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_16_nor_12_tmp, IsNaN_6U_10U_16_nor_12_itm,
          and_dcpl_547);
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_tmp,
          IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm, and_dcpl_547);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= 1'b0;
    end
    else if ( FpExpoWidthDec_6U_5U_10U_1U_1U_if_and_16_cse ) begin
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
          <= MUX_s_1_2_2(data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1,
          data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st,
          and_dcpl_547);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_mux1h_410_itm_4 <= 1'b0;
      data_truncate_nor_dfs_4 <= 1'b0;
      data_truncate_equal_tmp_4 <= 1'b0;
      data_truncate_nor_tmp_5 <= 1'b0;
      data_truncate_mux1h_320_itm_4 <= 1'b0;
      data_truncate_mux1h_404_itm_4 <= 1'b0;
      data_truncate_mux1h_326_itm_4 <= 1'b0;
      data_truncate_mux1h_398_itm_4 <= 1'b0;
      data_truncate_mux1h_332_itm_4 <= 1'b0;
      data_truncate_mux1h_392_itm_4 <= 1'b0;
      data_truncate_mux1h_338_itm_4 <= 1'b0;
      data_truncate_mux1h_386_itm_4 <= 1'b0;
      data_truncate_mux1h_344_itm_4 <= 1'b0;
      data_truncate_mux1h_380_itm_4 <= 1'b0;
      data_truncate_mux1h_350_itm_4 <= 1'b0;
      data_truncate_mux1h_374_itm_4 <= 1'b0;
      data_truncate_mux1h_356_itm_4 <= 1'b0;
      data_truncate_mux1h_368_itm_4 <= 1'b0;
      data_truncate_mux1h_362_itm_4 <= 1'b0;
    end
    else if ( data_truncate_and_cse ) begin
      data_truncate_mux1h_410_itm_4 <= data_truncate_mux1h_410_itm_3;
      data_truncate_nor_dfs_4 <= data_truncate_nor_dfs_3;
      data_truncate_equal_tmp_4 <= data_truncate_equal_tmp_3;
      data_truncate_nor_tmp_5 <= data_truncate_nor_tmp_4;
      data_truncate_mux1h_320_itm_4 <= data_truncate_mux1h_320_itm_3;
      data_truncate_mux1h_404_itm_4 <= data_truncate_mux1h_404_itm_3;
      data_truncate_mux1h_326_itm_4 <= data_truncate_mux1h_326_itm_3;
      data_truncate_mux1h_398_itm_4 <= data_truncate_mux1h_398_itm_3;
      data_truncate_mux1h_332_itm_4 <= data_truncate_mux1h_332_itm_3;
      data_truncate_mux1h_392_itm_4 <= data_truncate_mux1h_392_itm_3;
      data_truncate_mux1h_338_itm_4 <= data_truncate_mux1h_338_itm_3;
      data_truncate_mux1h_386_itm_4 <= data_truncate_mux1h_386_itm_3;
      data_truncate_mux1h_344_itm_4 <= data_truncate_mux1h_344_itm_3;
      data_truncate_mux1h_380_itm_4 <= data_truncate_mux1h_380_itm_3;
      data_truncate_mux1h_350_itm_4 <= data_truncate_mux1h_350_itm_3;
      data_truncate_mux1h_374_itm_4 <= data_truncate_mux1h_374_itm_3;
      data_truncate_mux1h_356_itm_4 <= data_truncate_mux1h_356_itm_3;
      data_truncate_mux1h_368_itm_4 <= data_truncate_mux1h_368_itm_3;
      data_truncate_mux1h_362_itm_4 <= data_truncate_mux1h_362_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_0_6_1_sva_10 <= 6'b0;
      o_data_data_15_13_10_sva_6 <= 4'b0;
      o_data_data_0_9_7_sva_6 <= 3'b0;
      o_data_data_15_9_7_sva_6 <= 3'b0;
      o_data_data_0_13_10_sva_6 <= 4'b0;
      o_data_data_15_6_1_sva_10 <= 6'b0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_1_6_1_sva_10 <= 6'b0;
      o_data_data_14_13_10_sva_6 <= 4'b0;
      o_data_data_1_9_7_sva_6 <= 3'b0;
      o_data_data_14_9_7_sva_6 <= 3'b0;
      o_data_data_1_13_10_sva_6 <= 4'b0;
      o_data_data_14_6_1_sva_10 <= 6'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_2_6_1_sva_10 <= 6'b0;
      o_data_data_13_13_10_sva_6 <= 4'b0;
      o_data_data_2_9_7_sva_6 <= 3'b0;
      o_data_data_13_9_7_sva_6 <= 3'b0;
      o_data_data_2_13_10_sva_6 <= 4'b0;
      o_data_data_13_6_1_sva_10 <= 6'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_3_6_1_sva_10 <= 6'b0;
      o_data_data_12_13_10_sva_6 <= 4'b0;
      o_data_data_3_9_7_sva_6 <= 3'b0;
      o_data_data_12_9_7_sva_6 <= 3'b0;
      o_data_data_3_13_10_sva_6 <= 4'b0;
      o_data_data_12_6_1_sva_10 <= 6'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_4_6_1_sva_10 <= 6'b0;
      o_data_data_11_13_10_sva_6 <= 4'b0;
      o_data_data_4_9_7_sva_6 <= 3'b0;
      o_data_data_11_9_7_sva_6 <= 3'b0;
      o_data_data_4_13_10_sva_6 <= 4'b0;
      o_data_data_11_6_1_sva_10 <= 6'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_5_6_1_sva_10 <= 6'b0;
      o_data_data_10_13_10_sva_6 <= 4'b0;
      o_data_data_5_9_7_sva_6 <= 3'b0;
      o_data_data_10_9_7_sva_6 <= 3'b0;
      o_data_data_5_13_10_sva_6 <= 4'b0;
      o_data_data_10_6_1_sva_10 <= 6'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_6_6_1_sva_10 <= 6'b0;
      o_data_data_9_13_10_sva_6 <= 4'b0;
      o_data_data_6_9_7_sva_6 <= 3'b0;
      o_data_data_9_9_7_sva_6 <= 3'b0;
      o_data_data_6_13_10_sva_6 <= 4'b0;
      o_data_data_9_6_1_sva_10 <= 6'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      o_data_data_7_6_1_sva_10 <= 6'b0;
      o_data_data_8_13_10_sva_6 <= 4'b0;
      o_data_data_7_9_7_sva_6 <= 3'b0;
      o_data_data_8_9_7_sva_6 <= 3'b0;
      o_data_data_7_13_10_sva_6 <= 4'b0;
      o_data_data_8_6_1_sva_10 <= 6'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= 1'b0;
    end
    else if ( IntShiftRight_18U_2U_16U_obits_fixed_and_16_cse ) begin
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_0_6_1_sva_10 <= o_data_data_0_6_1_sva_9;
      o_data_data_15_13_10_sva_6 <= o_data_data_15_13_10_sva_5;
      o_data_data_0_9_7_sva_6 <= o_data_data_0_9_7_sva_5;
      o_data_data_15_9_7_sva_6 <= o_data_data_15_9_7_sva_5;
      o_data_data_0_13_10_sva_6 <= o_data_data_0_13_10_sva_5;
      o_data_data_15_6_1_sva_10 <= o_data_data_15_6_1_sva_9;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_1_6_1_sva_10 <= o_data_data_1_6_1_sva_9;
      o_data_data_14_13_10_sva_6 <= o_data_data_14_13_10_sva_5;
      o_data_data_1_9_7_sva_6 <= o_data_data_1_9_7_sva_5;
      o_data_data_14_9_7_sva_6 <= o_data_data_14_9_7_sva_5;
      o_data_data_1_13_10_sva_6 <= o_data_data_1_13_10_sva_5;
      o_data_data_14_6_1_sva_10 <= o_data_data_14_6_1_sva_9;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_2_6_1_sva_10 <= o_data_data_2_6_1_sva_9;
      o_data_data_13_13_10_sva_6 <= o_data_data_13_13_10_sva_5;
      o_data_data_2_9_7_sva_6 <= o_data_data_2_9_7_sva_5;
      o_data_data_13_9_7_sva_6 <= o_data_data_13_9_7_sva_5;
      o_data_data_2_13_10_sva_6 <= o_data_data_2_13_10_sva_5;
      o_data_data_13_6_1_sva_10 <= o_data_data_13_6_1_sva_9;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_3_6_1_sva_10 <= o_data_data_3_6_1_sva_9;
      o_data_data_12_13_10_sva_6 <= o_data_data_12_13_10_sva_5;
      o_data_data_3_9_7_sva_6 <= o_data_data_3_9_7_sva_5;
      o_data_data_12_9_7_sva_6 <= o_data_data_12_9_7_sva_5;
      o_data_data_3_13_10_sva_6 <= o_data_data_3_13_10_sva_5;
      o_data_data_12_6_1_sva_10 <= o_data_data_12_6_1_sva_9;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_4_6_1_sva_10 <= o_data_data_4_6_1_sva_9;
      o_data_data_11_13_10_sva_6 <= o_data_data_11_13_10_sva_5;
      o_data_data_4_9_7_sva_6 <= o_data_data_4_9_7_sva_5;
      o_data_data_11_9_7_sva_6 <= o_data_data_11_9_7_sva_5;
      o_data_data_4_13_10_sva_6 <= o_data_data_4_13_10_sva_5;
      o_data_data_11_6_1_sva_10 <= o_data_data_11_6_1_sva_9;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_5_6_1_sva_10 <= o_data_data_5_6_1_sva_9;
      o_data_data_10_13_10_sva_6 <= o_data_data_10_13_10_sva_5;
      o_data_data_5_9_7_sva_6 <= o_data_data_5_9_7_sva_5;
      o_data_data_10_9_7_sva_6 <= o_data_data_10_9_7_sva_5;
      o_data_data_5_13_10_sva_6 <= o_data_data_5_13_10_sva_5;
      o_data_data_10_6_1_sva_10 <= o_data_data_10_6_1_sva_9;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_6_6_1_sva_10 <= o_data_data_6_6_1_sva_9;
      o_data_data_9_13_10_sva_6 <= o_data_data_9_13_10_sva_5;
      o_data_data_6_9_7_sva_6 <= o_data_data_6_9_7_sva_5;
      o_data_data_9_9_7_sva_6 <= o_data_data_9_9_7_sva_5;
      o_data_data_6_13_10_sva_6 <= o_data_data_6_13_10_sva_5;
      o_data_data_9_6_1_sva_10 <= o_data_data_9_6_1_sva_9;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      o_data_data_7_6_1_sva_10 <= o_data_data_7_6_1_sva_9;
      o_data_data_8_13_10_sva_6 <= o_data_data_8_13_10_sva_5;
      o_data_data_7_9_7_sva_6 <= o_data_data_7_9_7_sva_5;
      o_data_data_8_9_7_sva_6 <= o_data_data_8_9_7_sva_5;
      o_data_data_7_13_10_sva_6 <= o_data_data_7_13_10_sva_5;
      o_data_data_8_6_1_sva_10 <= o_data_data_8_6_1_sva_9;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_4
          <= data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_4
          <= data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_0_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_15_6_1_sva_8 <= 6'b0;
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_1_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_14_6_1_sva_8 <= 6'b0;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_2_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_13_6_1_sva_8 <= 6'b0;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_3_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_12_6_1_sva_8 <= 6'b0;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_4_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_11_6_1_sva_8 <= 6'b0;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_5_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_10_6_1_sva_8 <= 6'b0;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_6_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_9_6_1_sva_8 <= 6'b0;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= 1'b0;
      o_data_data_7_6_1_sva_8 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= 1'b0;
      o_data_data_8_6_1_sva_8 <= 6'b0;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= 1'b0;
    end
    else if ( IntShiftRight_18U_2U_8U_obits_fixed_and_16_cse ) begin
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_0_6_1_sva_8 <= o_data_data_0_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_15_6_1_sva_8 <= o_data_data_15_6_1_sva_7;
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_1_6_1_sva_8 <= o_data_data_1_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_14_6_1_sva_8 <= o_data_data_14_6_1_sva_7;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_2_6_1_sva_8 <= o_data_data_2_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_13_6_1_sva_8 <= o_data_data_13_6_1_sva_7;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_3_6_1_sva_8 <= o_data_data_3_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_12_6_1_sva_8 <= o_data_data_12_6_1_sva_7;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_4_6_1_sva_8 <= o_data_data_4_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_11_6_1_sva_8 <= o_data_data_11_6_1_sva_7;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_5_6_1_sva_8 <= o_data_data_5_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_10_6_1_sva_8 <= o_data_data_10_6_1_sva_7;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_6_6_1_sva_8 <= o_data_data_6_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_9_6_1_sva_8 <= o_data_data_9_6_1_sva_7;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_7_6_1_sva_8 <= o_data_data_7_6_1_sva_7;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_5_itm_4
          <= IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3;
      o_data_data_8_6_1_sva_8 <= o_data_data_8_6_1_sva_7;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_4
          <= data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_mant_3_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_211_nl) ) begin
      FpAdd_6U_10U_7_o_mant_3_lpi_2 <= FpAdd_6U_10U_7_o_mant_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_mant_2_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_215_nl) ) begin
      FpAdd_6U_10U_7_o_mant_2_lpi_2 <= FpAdd_6U_10U_7_o_mant_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_mant_1_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_218_nl) ) begin
      FpAdd_6U_10U_7_o_mant_1_lpi_2 <= FpAdd_6U_10U_7_o_mant_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_expo_3_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_227_nl) ) begin
      FpAdd_6U_10U_7_o_expo_3_lpi_2 <= FpAdd_6U_10U_7_o_expo_3_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_expo_2_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_236_nl) ) begin
      FpAdd_6U_10U_7_o_expo_2_lpi_2 <= FpAdd_6U_10U_7_o_expo_2_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_expo_1_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_245_nl) ) begin
      FpAdd_6U_10U_7_o_expo_1_lpi_2 <= FpAdd_6U_10U_7_o_expo_1_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_mant_3_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_249_nl) ) begin
      FpAdd_6U_10U_6_o_mant_3_lpi_2 <= FpAdd_6U_10U_6_o_mant_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_mant_2_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_253_nl) ) begin
      FpAdd_6U_10U_6_o_mant_2_lpi_2 <= FpAdd_6U_10U_6_o_mant_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_mant_1_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_257_nl) ) begin
      FpAdd_6U_10U_6_o_mant_1_lpi_2 <= FpAdd_6U_10U_6_o_mant_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_expo_3_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_266_nl) ) begin
      FpAdd_6U_10U_6_o_expo_3_lpi_2 <= FpAdd_6U_10U_6_o_expo_3_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_expo_2_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_275_nl) ) begin
      FpAdd_6U_10U_6_o_expo_2_lpi_2 <= FpAdd_6U_10U_6_o_expo_2_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_expo_1_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_284_nl) ) begin
      FpAdd_6U_10U_6_o_expo_1_lpi_2 <= FpAdd_6U_10U_6_o_expo_1_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_mant_3_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_289_nl) ) begin
      FpAdd_6U_10U_5_o_mant_3_lpi_2 <= FpAdd_6U_10U_5_o_mant_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_mant_2_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_295_nl) ) begin
      FpAdd_6U_10U_5_o_mant_2_lpi_2 <= FpAdd_6U_10U_5_o_mant_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_mant_1_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_298_nl) ) begin
      FpAdd_6U_10U_5_o_mant_1_lpi_2 <= FpAdd_6U_10U_5_o_mant_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_expo_3_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_307_nl) ) begin
      FpAdd_6U_10U_5_o_expo_3_lpi_2 <= FpAdd_6U_10U_5_o_expo_3_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_expo_2_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_316_nl) ) begin
      FpAdd_6U_10U_5_o_expo_2_lpi_2 <= FpAdd_6U_10U_5_o_expo_2_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_expo_1_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_325_nl) ) begin
      FpAdd_6U_10U_5_o_expo_1_lpi_2 <= FpAdd_6U_10U_5_o_expo_1_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_mant_3_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_328_nl) ) begin
      FpAdd_6U_10U_4_o_mant_3_lpi_2 <= FpAdd_6U_10U_4_o_mant_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_mant_2_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_334_nl) ) begin
      FpAdd_6U_10U_4_o_mant_2_lpi_2 <= FpAdd_6U_10U_4_o_mant_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_mant_1_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_339_nl) ) begin
      FpAdd_6U_10U_4_o_mant_1_lpi_2 <= FpAdd_6U_10U_4_o_mant_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_expo_3_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_348_nl) ) begin
      FpAdd_6U_10U_4_o_expo_3_lpi_2 <= FpAdd_6U_10U_4_o_expo_3_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_expo_2_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_354_nl) ) begin
      FpAdd_6U_10U_4_o_expo_2_lpi_2 <= FpAdd_6U_10U_4_o_expo_2_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_expo_1_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_363_nl) ) begin
      FpAdd_6U_10U_4_o_expo_1_lpi_2 <= FpAdd_6U_10U_4_o_expo_1_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_mant_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_370_nl) ) begin
      FpAdd_6U_10U_7_o_mant_lpi_2 <= FpAdd_6U_10U_7_o_mant_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_expo_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_379_nl) ) begin
      FpAdd_6U_10U_7_o_expo_lpi_2 <= FpAdd_6U_10U_7_o_expo_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_mant_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_383_nl) ) begin
      FpAdd_6U_10U_6_o_mant_lpi_2 <= FpAdd_6U_10U_6_o_mant_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_6_o_expo_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_392_nl) ) begin
      FpAdd_6U_10U_6_o_expo_lpi_2 <= FpAdd_6U_10U_6_o_expo_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_mant_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_396_nl) ) begin
      FpAdd_6U_10U_5_o_mant_lpi_2 <= FpAdd_6U_10U_5_o_mant_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_5_o_expo_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_405_nl) ) begin
      FpAdd_6U_10U_5_o_expo_lpi_2 <= FpAdd_6U_10U_5_o_expo_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_mant_lpi_2 <= 10'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_412_nl) ) begin
      FpAdd_6U_10U_4_o_mant_lpi_2 <= FpAdd_6U_10U_4_o_mant_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_4_o_expo_lpi_2 <= 6'b0;
    end
    else if ( core_wen & (~ or_dcpl_296) & (mux_421_nl) ) begin
      FpAdd_6U_10U_4_o_expo_lpi_2 <= FpAdd_6U_10U_4_o_expo_lpi_1_dfm_8_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm <= 1'b0;
      IsNaN_6U_10U_16_nor_15_itm <= 1'b0;
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm <= 1'b0;
      IsNaN_6U_10U_16_nor_12_itm <= 1'b0;
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= 1'b0;
    end
    else if ( IsNaN_6U_10U_16_and_cse ) begin
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_tmp;
      IsNaN_6U_10U_16_nor_15_itm <= IsNaN_6U_10U_16_nor_15_tmp;
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm <= IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_tmp;
      IsNaN_6U_10U_16_nor_12_itm <= IsNaN_6U_10U_16_nor_12_tmp;
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
          <= data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st <= 1'b0;
      IsNaN_6U_10U_14_land_lpi_1_dfm_st <= 1'b0;
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= 1'b0;
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= 1'b0;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_st <= 1'b0;
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= 1'b0;
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= 1'b0;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_st <= 1'b0;
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= 1'b0;
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= 1'b0;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_st <= 1'b0;
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= 1'b0;
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= 1'b0;
      IsNaN_6U_10U_12_land_lpi_1_dfm_st <= 1'b0;
      o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= 1'b0;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st <= 1'b0;
      o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= 1'b0;
      o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= 1'b0;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st <= 1'b0;
      o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= 1'b0;
      o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= 1'b0;
      o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= 1'b0;
      o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= 1'b0;
      o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= 1'b0;
    end
    else if ( IsNaN_6U_10U_12_aelse_and_cse ) begin
      IsNaN_6U_10U_12_land_2_lpi_1_dfm_st <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp;
      IsNaN_6U_10U_14_land_lpi_1_dfm_st <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp;
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
      o_col3_4_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= o_col1_4_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
      IsNaN_6U_10U_14_land_3_lpi_1_dfm_st <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp;
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
      o_col3_3_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= o_col1_3_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
      IsNaN_6U_10U_14_land_2_lpi_1_dfm_st <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp;
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
      o_col3_2_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= o_col1_2_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
      IsNaN_6U_10U_14_land_1_lpi_1_dfm_st <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp;
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm <= o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_15_or_itm_mx0w0;
      o_col3_1_FpAdd_6U_10U_7_IsZero_6U_10U_14_or_itm <= o_col1_1_FpAdd_6U_10U_5_IsZero_6U_10U_10_or_itm_mx0w0;
      IsNaN_6U_10U_12_land_lpi_1_dfm_st <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp;
      o_col2_4_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
      IsNaN_6U_10U_12_land_3_lpi_1_dfm_st <= IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp;
      o_col2_3_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
      o_col2_2_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
      IsNaN_6U_10U_12_land_1_lpi_1_dfm_st <= IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp;
      o_col2_1_FpAdd_6U_10U_6_IsZero_6U_10U_12_or_itm <= o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_9_or_itm_mx0w0;
      o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= o_col0_4_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
      o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= o_col0_3_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
      o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= o_col0_2_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
      o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm <= o_col0_1_FpAdd_6U_10U_4_IsZero_6U_10U_8_or_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2 <= 10'b0;
    end
    else if ( core_wen & ((and_tmp_56 & and_dcpl_88 & reg_IsNaN_6U_10U_6_land_lpi_1_dfm_st_1_cse)
        | FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx0c1) ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_3_FpAdd_6U_10U_3_or_11_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_8_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2 <= 10'b0;
    end
    else if ( core_wen & ((and_tmp_56 & and_dcpl_88 & IsNaN_6U_10U_4_land_lpi_1_dfm_st_2)
        | FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx0c1) ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_2_FpAdd_6U_10U_2_or_11_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_8_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2 <= 10'b0;
    end
    else if ( core_wen & ((and_tmp_56 & and_dcpl_88 & IsNaN_6U_10U_2_land_lpi_1_dfm_st_2)
        | FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx0c1) ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_11_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_8_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_2 <= 10'b0;
    end
    else if ( core_wen & ((and_tmp_56 & and_dcpl_88 & reg_IsNaN_6U_10U_land_lpi_1_dfm_st_1_cse)
        | FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0c1) ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_2 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7,
          FpAdd_6U_10U_FpAdd_6U_10U_or_11_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_932_rgt | and_935_rgt | and_938_rgt | and_941_rgt)
        & mux_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[137:128]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          (chn_data_in_rsci_d_mxwt[9:0]), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w4,
          {and_932_rgt , and_935_rgt , and_938_rgt , and_941_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_9_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_5 <= MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3, and_dcpl_658);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2, and_dcpl_658);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_IsNaN_6U_10U_and_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm <= IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_946_rgt | and_949_rgt | and_952_rgt | and_955_rgt)
        & (mux_2_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[153:144]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          (chn_data_in_rsci_d_mxwt[25:16]), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_2_mx0w4,
          {and_946_rgt , and_949_rgt , and_952_rgt , and_955_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_11_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_5 <= MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3, and_dcpl_672);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2, and_dcpl_672);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm <= IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_960_rgt | and_963_rgt | and_966_rgt | and_969_rgt)
        & mux_9_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[169:160]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          (chn_data_in_rsci_d_mxwt[41:32]), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w4,
          {and_960_rgt , and_963_rgt , and_966_rgt , and_969_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_5 <= MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3, and_dcpl_686);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2, and_dcpl_686);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | (cfg_precision[0]) | IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp
        | (~ chn_data_in_rsci_bawt) | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm <= IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_974_rgt | and_977_rgt | and_980_rgt | and_983_rgt)
        & mux_13_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[73:64]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          (chn_data_in_rsci_d_mxwt[137:128]), FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          {and_974_rgt , and_977_rgt , and_980_rgt , and_983_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_14_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_687) | and_985_rgt) & mux_13_cse
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, and_985_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_988_rgt | and_991_rgt | and_994_rgt | and_997_rgt)
        & mux_16_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[89:80]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          (chn_data_in_rsci_d_mxwt[153:144]), FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          {and_988_rgt , and_991_rgt , and_994_rgt , and_997_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_17_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_701) | and_999_rgt) & mux_16_cse
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, and_999_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_2_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1002_rgt | and_1005_rgt | and_1008_rgt | and_1011_rgt)
        & (mux_21_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[105:96]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          (chn_data_in_rsci_d_mxwt[169:160]), FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          {and_1002_rgt , and_1005_rgt , and_1008_rgt , and_1011_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_22_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_715) | and_1013_rgt) & (mux_23_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, and_1013_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_4_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1016_rgt | and_1019_rgt | and_1022_rgt | and_1025_rgt)
        & mux_27_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_1_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[137:128]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_mx0w1,
          (chn_data_in_rsci_d_mxwt[73:64]), FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          {and_1016_rgt , and_1019_rgt , and_1022_rgt , and_1025_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_6 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_9_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, and_dcpl_742);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]), and_dcpl_742);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          and_dcpl_742);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1030_rgt | and_1033_rgt | and_1036_rgt | and_1039_rgt)
        & mux_29_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_2_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[153:144]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_2_mx0w1,
          (chn_data_in_rsci_d_mxwt[89:80]), FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          {and_1030_rgt , and_1033_rgt , and_1036_rgt , and_1039_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_6 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_10_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, and_dcpl_756);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]), and_dcpl_756);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          and_dcpl_756);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1044_rgt | and_1047_rgt | and_1050_rgt | and_1053_rgt)
        & mux_31_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_3_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[169:160]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_4_mx0w1,
          (chn_data_in_rsci_d_mxwt[105:96]), FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          {and_1044_rgt , and_1047_rgt , and_1050_rgt , and_1053_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_6 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_11_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, and_dcpl_770);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]), and_dcpl_770);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          and_dcpl_770);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1058_rgt | and_1061_rgt | and_1064_rgt | and_1067_rgt)
        & (mux_36_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_1_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[73:64]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_mx0w1,
          (chn_data_in_rsci_d_mxwt[201:192]), FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_mx0w4,
          {and_1058_rgt , and_1061_rgt , and_1064_rgt , and_1067_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_771) | and_1069_rgt) & (mux_37_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2, and_1069_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (~ (mux_39_nl)) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm <= IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1072_rgt | and_1075_rgt | and_1078_rgt | and_1081_rgt)
        & mux_40_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_2_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[89:80]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_2_mx0w1,
          (chn_data_in_rsci_d_mxwt[217:208]), FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_2_mx0w4,
          {and_1072_rgt , and_1075_rgt , and_1078_rgt , and_1081_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_785) | and_1083_rgt) & mux_40_cse
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2, and_1083_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_42_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm <= IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1086_rgt | and_1089_rgt | and_1092_rgt | and_1095_rgt)
        & (mux_43_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_3_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[105:96]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_4_mx0w1,
          (chn_data_in_rsci_d_mxwt[233:224]), FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_4_mx0w4,
          {and_1086_rgt , and_1089_rgt , and_1092_rgt , and_1095_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_799) | and_1097_rgt) & (mux_44_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2, and_1097_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_45_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm <= IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_6_land_lpi_1_dfm_st <= 1'b0;
      m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_6_land_3_lpi_1_dfm <= 1'b0;
      m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_6_land_2_lpi_1_dfm <= 1'b0;
      m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_6_land_1_lpi_1_dfm <= 1'b0;
      m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_4_land_lpi_1_dfm_st <= 1'b0;
      m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_4_land_3_lpi_1_dfm <= 1'b0;
      m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_4_land_2_lpi_1_dfm <= 1'b0;
      m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_4_land_1_lpi_1_dfm <= 1'b0;
      m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st <= 1'b0;
      m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm <= 1'b0;
      m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm <= 1'b0;
      m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm <= 1'b0;
      m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_st <= 1'b0;
      m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_land_3_lpi_1_dfm <= 1'b0;
      m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_land_2_lpi_1_dfm <= 1'b0;
      m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= 1'b0;
      IsNaN_6U_10U_land_1_lpi_1_dfm <= 1'b0;
      m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= 1'b0;
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= 1'b0;
      o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= 1'b0;
      o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= 1'b0;
      o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= 1'b0;
      o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= 1'b0;
      o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= 1'b0;
      o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= 1'b0;
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= 1'b0;
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= 1'b0;
      o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= 1'b0;
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= 1'b0;
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= 1'b0;
      o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= 1'b0;
      o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= 1'b0;
      o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= 1'b0;
      o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= 1'b0;
    end
    else if ( IsNaN_6U_10U_6_aelse_and_cse ) begin
      IsNaN_6U_10U_6_land_lpi_1_dfm_st <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
      m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= m_row3_4_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_6_land_3_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
      m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= m_row3_3_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_6_land_2_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp;
      m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= m_row3_2_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_6_land_1_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
      m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_st
          <= m_row3_1_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_FpAdd_6U_10U_3_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_4_land_lpi_1_dfm_st <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
      m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= m_row2_4_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_4_land_3_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp;
      m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= m_row2_3_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_4_land_2_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp;
      m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= m_row2_2_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_4_land_1_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp;
      m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_st
          <= m_row2_1_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_FpAdd_6U_10U_2_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st <= IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp;
      m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= m_row1_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm <= IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp;
      m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= m_row1_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm <= IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp;
      m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= m_row1_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm <= IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp;
      m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st
          <= m_row1_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
      IsNaN_6U_10U_land_lpi_1_dfm_st <= IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp;
      m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= m_row0_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_land_3_lpi_1_dfm <= IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp;
      m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= m_row0_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_land_2_lpi_1_dfm <= IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp;
      m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= m_row0_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
      IsNaN_6U_10U_land_1_lpi_1_dfm <= IsNaN_6U_10U_IsNaN_6U_10U_and_tmp;
      m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_st
          <= m_row0_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xor_svs_mx0w0;
      o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= o_col3_4_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
      o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= o_col3_3_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
      o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= o_col3_2_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
      o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_st
          <= o_col3_1_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_FpAdd_6U_10U_7_is_addition_xor_svs_mx0w0;
      o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= o_col2_4_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
      o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= o_col2_3_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
      o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= o_col2_2_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
      o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_st
          <= o_col2_1_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_FpAdd_6U_10U_6_is_addition_xor_svs_mx0w0;
      o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= o_col1_4_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
      o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= o_col1_3_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
      o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= o_col1_2_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
      o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_st
          <= o_col1_1_FpAdd_6U_10U_5_is_addition_FpAdd_6U_10U_5_is_addition_xnor_svs_mx0w0;
      o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= o_col0_4_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
      o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= o_col0_3_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
      o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= o_col0_2_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
      o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_st
          <= o_col0_1_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_FpAdd_6U_10U_4_is_addition_xor_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_b_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_b_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_3_a_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_b_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_2_a_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_1_a_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_b_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_a_int_mant_p1_sva <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_b_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_a_int_mant_p1_3_sva <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_b_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_a_int_mant_p1_2_sva <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_b_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_a_int_mant_p1_1_sva <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_4_cse ) begin
      FpAdd_6U_10U_3_b_int_mant_p1_sva <= FpAdd_6U_10U_3_b_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_3_a_int_mant_p1_sva <= FpAdd_6U_10U_3_a_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_3_is_a_greater_lor_lpi_1_dfm_1 <= FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp;
      FpAdd_6U_10U_3_b_int_mant_p1_3_sva <= FpAdd_6U_10U_3_b_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_3_a_int_mant_p1_3_sva <= FpAdd_6U_10U_3_a_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_3_is_a_greater_lor_3_lpi_1_dfm_1 <= FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp;
      FpAdd_6U_10U_3_b_int_mant_p1_2_sva <= FpAdd_6U_10U_3_b_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_3_a_int_mant_p1_2_sva <= FpAdd_6U_10U_3_a_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_3_is_a_greater_lor_2_lpi_1_dfm_1 <= FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp;
      FpAdd_6U_10U_3_b_int_mant_p1_1_sva <= FpAdd_6U_10U_3_b_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_3_a_int_mant_p1_1_sva <= FpAdd_6U_10U_3_a_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_3_is_a_greater_lor_1_lpi_1_dfm_1 <= FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp;
      FpAdd_6U_10U_2_b_int_mant_p1_sva <= FpAdd_6U_10U_2_b_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_2_a_int_mant_p1_sva <= FpAdd_6U_10U_2_a_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_2_is_a_greater_lor_lpi_1_dfm_1 <= FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp;
      FpAdd_6U_10U_2_b_int_mant_p1_3_sva <= FpAdd_6U_10U_2_b_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_2_a_int_mant_p1_3_sva <= FpAdd_6U_10U_2_a_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_2_is_a_greater_lor_3_lpi_1_dfm_1 <= FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp;
      FpAdd_6U_10U_2_b_int_mant_p1_2_sva <= FpAdd_6U_10U_2_b_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_2_a_int_mant_p1_2_sva <= FpAdd_6U_10U_2_a_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_2_is_a_greater_lor_2_lpi_1_dfm_1 <= FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp;
      FpAdd_6U_10U_2_b_int_mant_p1_1_sva <= FpAdd_6U_10U_2_b_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_2_a_int_mant_p1_1_sva <= FpAdd_6U_10U_2_a_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_2_is_a_greater_lor_1_lpi_1_dfm_1 <= FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp;
      FpAdd_6U_10U_1_b_int_mant_p1_sva <= FpAdd_6U_10U_1_b_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_1_a_int_mant_p1_sva <= FpAdd_6U_10U_1_a_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1 <= FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp;
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva <= FpAdd_6U_10U_1_b_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_1_a_int_mant_p1_3_sva <= FpAdd_6U_10U_1_a_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1 <= FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp;
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva <= FpAdd_6U_10U_1_b_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_1_a_int_mant_p1_2_sva <= FpAdd_6U_10U_1_a_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1 <= FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp;
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva <= FpAdd_6U_10U_1_b_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_1_a_int_mant_p1_1_sva <= FpAdd_6U_10U_1_a_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1 <= FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp;
      FpAdd_6U_10U_b_int_mant_p1_sva <= FpAdd_6U_10U_b_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_a_int_mant_p1_sva <= FpAdd_6U_10U_a_int_mant_p1_sva_mx0w0;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1 <= FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp;
      FpAdd_6U_10U_b_int_mant_p1_3_sva <= FpAdd_6U_10U_b_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_a_int_mant_p1_3_sva <= FpAdd_6U_10U_a_int_mant_p1_3_sva_mx0w0;
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1 <= FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp;
      FpAdd_6U_10U_b_int_mant_p1_2_sva <= FpAdd_6U_10U_b_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_a_int_mant_p1_2_sva <= FpAdd_6U_10U_a_int_mant_p1_2_sva_mx0w0;
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1 <= FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp;
      FpAdd_6U_10U_b_int_mant_p1_1_sva <= FpAdd_6U_10U_b_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_a_int_mant_p1_1_sva <= FpAdd_6U_10U_a_int_mant_p1_1_sva_mx0w0;
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1 <= FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1769_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp)
        | FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_and_29_cse ) begin
      FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4[1]), and_1771_cse);
      FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4[0]), and_1771_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_12_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_3_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1801_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp)
        | FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_3_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_and_32_cse ) begin
      FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4[1]), and_1803_cse);
      FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4[0]), and_1803_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_14_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_2_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1833_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp)
        | FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_2_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_and_35_cse ) begin
      FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4[1]), and_1835_cse);
      FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4[0]), and_1835_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_16_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_1_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1865_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp)
        | FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_1_lpi_1_dfm_3_mx0w2, FpAdd_6U_10U_3_qr_3_0_1_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_and_38_cse ) begin
      FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4[1]), and_1867_cse);
      FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4[0]), and_1867_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1895_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp)
        | FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_2_and_29_cse ) begin
      FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]), and_1897_cse);
      FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          and_1897_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1927_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp)
        | FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_2_and_32_cse ) begin
      FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]), and_1929_cse);
      FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          and_1929_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1959_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp)
        | FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_2_and_35_cse ) begin
      FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]), and_1961_cse);
      FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          and_1961_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_1991_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp)
        | FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_2_qr_3_0_1_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_2_and_38_cse ) begin
      FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]), and_1993_cse);
      FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          and_1993_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2021_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp)
        | FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_and_29_cse ) begin
      FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]), and_2023_cse);
      FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          and_2023_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2053_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_2_tmp)
        | FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_and_32_cse ) begin
      FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]), and_2055_cse);
      FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          and_2055_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2085_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_1_tmp)
        | FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_and_35_cse ) begin
      FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]), and_2087_cse);
      FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          and_2087_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2117_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp)
        | FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_1_qr_3_0_1_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_and_38_cse ) begin
      FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]), and_2119_cse);
      FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          and_2119_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2147_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp)
        | FpAdd_6U_10U_qr_3_0_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_qr_3_0_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_5_4_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_qr_5_4_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_29_cse ) begin
      FpAdd_6U_10U_qr_5_4_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]), and_2149_cse);
      FpAdd_6U_10U_qr_5_4_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[0]), and_2149_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2179_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp)
        | FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_3_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_32_cse ) begin
      FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]), and_2181_cse);
      FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[0]), and_2181_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2211_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp)
        | FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_2_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_35_cse ) begin
      FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]), and_2213_cse);
      FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[0]), and_2213_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm <= 4'b0;
    end
    else if ( core_wen & (and_2243_cse | (and_dcpl_817 & and_dcpl_57 & FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp)
        | FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_mx0c1) ) begin
      FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w2,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_1_lpi_1_dfm_3_mx0w0, FpAdd_6U_10U_qr_3_0_1_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_1 <= 1'b0;
      FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_0 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_38_cse ) begin
      FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]), and_2245_cse);
      FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_0 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[0]), and_2245_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_1268_rgt | and_1271_rgt | and_dcpl_78 | and_1280_rgt
        | and_1283_rgt) & (mux_434_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[185:176]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[57:48]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_6_mx0w4,
          {and_1268_rgt , and_1271_rgt , and_dcpl_78 , and_1280_rgt , and_1283_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_999 | and_1285_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp,
          IsNaN_6U_10U_1_land_lpi_1_dfm, and_1285_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1002 | and_1288_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp,
          IsNaN_6U_10U_3_land_lpi_1_dfm, and_1288_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1005 | and_1291_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp,
          IsNaN_6U_10U_5_land_lpi_1_dfm, and_1291_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1008 | and_1294_rgt) & mux_tmp_49 ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp,
          IsNaN_6U_10U_7_land_lpi_1_dfm, and_1294_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_1303_rgt | and_1306_rgt | and_dcpl_78 | and_1314_rgt
        | and_1317_rgt) & (mux_440_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[121:112]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[249:240]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_6_mx0w4,
          {and_1303_rgt , and_1306_rgt , and_dcpl_78 , and_1314_rgt , and_1317_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_3_mx0[1]),
          {and_dcpl_1033 , and_dcpl_1034 , and_dcpl_1035});
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_0_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_3_mx0[0]),
          {and_dcpl_1033 , and_dcpl_1034 , and_dcpl_1035});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_1033 | and_dcpl_78 | and_dcpl_1008) & mux_tmp_443
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2,
          {and_dcpl_1033 , and_dcpl_78 , and_dcpl_1008});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_1323_rgt | and_1325_rgt | and_dcpl_78 | and_1327_rgt
        | and_1329_rgt) & (mux_446_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[185:176]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[121:112]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          {and_1323_rgt , and_1325_rgt , and_dcpl_78 , and_1327_rgt , and_1329_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_7 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_1_1, (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          {and_dcpl_1045 , and_dcpl_78 , and_dcpl_1005});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          {and_dcpl_1045 , and_dcpl_78 , and_dcpl_1005});
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          {and_dcpl_1045 , and_dcpl_78 , and_dcpl_1005});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (and_1333_rgt | and_1335_rgt | and_dcpl_78 | and_1337_rgt
        | and_1339_rgt) & (mux_453_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_7 <= MUX1HOT_v_10_5_2((chn_data_in_rsci_d_mxwt[121:112]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_6, (chn_data_in_rsci_d_mxwt[185:176]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          {and_1333_rgt , and_1335_rgt , and_dcpl_78 , and_1337_rgt , and_1339_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_1_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]), FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1_1,
          {and_dcpl_1055 , and_dcpl_1002 , and_dcpl_1056});
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5_0_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_mx0[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_1, {and_dcpl_1055
          , and_dcpl_1002 , and_dcpl_1056});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_1342_rgt | and_dcpl_78 | and_dcpl_1002) & mux_tmp_457
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          {and_1342_rgt , and_dcpl_78 , and_dcpl_1002});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_mx0[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_mx0[1]), and_dcpl_1059);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5_0_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_mx0[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_mx0[0]), and_dcpl_1059);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_7 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_999 | and_dcpl_78 | and_1345_rgt) & mux_tmp_460
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_7 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_6, FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2,
          {and_dcpl_999 , and_dcpl_78 , and_1345_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      o_data_data_15_6_1_sva_7 <= 6'b0;
      o_data_data_14_6_1_sva_7 <= 6'b0;
      o_data_data_13_6_1_sva_7 <= 6'b0;
      o_data_data_12_6_1_sva_7 <= 6'b0;
      o_data_data_11_6_1_sva_7 <= 6'b0;
      o_data_data_10_6_1_sva_7 <= 6'b0;
      o_data_data_9_6_1_sva_7 <= 6'b0;
      o_data_data_8_6_1_sva_7 <= 6'b0;
      o_data_data_7_6_1_sva_7 <= 6'b0;
      o_data_data_6_6_1_sva_7 <= 6'b0;
      o_data_data_5_6_1_sva_7 <= 6'b0;
      o_data_data_4_6_1_sva_7 <= 6'b0;
      o_data_data_3_6_1_sva_7 <= 6'b0;
      o_data_data_2_6_1_sva_7 <= 6'b0;
      o_data_data_1_6_1_sva_7 <= 6'b0;
      o_data_data_0_6_1_sva_7 <= 6'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= 1'b0;
    end
    else if ( o_data_data_and_64_cse ) begin
      o_data_data_15_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_sva));
      o_data_data_14_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_15_sva));
      o_data_data_13_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_14_sva));
      o_data_data_12_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_13_sva));
      o_data_data_11_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_12_sva));
      o_data_data_10_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_11_sva));
      o_data_data_9_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_10_sva));
      o_data_data_8_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_9_sva));
      o_data_data_7_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_8_sva));
      o_data_data_6_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_7_sva));
      o_data_data_5_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_6_sva));
      o_data_data_4_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_5_sva));
      o_data_data_3_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_4_sva));
      o_data_data_2_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_3_sva));
      o_data_data_1_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_2_sva));
      o_data_data_0_6_1_sva_7 <= ~(MUX_v_6_2_2((data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl),
          6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_1_sva));
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out[17];
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_1[17];
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_1[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_15_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_15_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_2[17];
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_2[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_14_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_14_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_3[17];
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_3[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_13_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_13_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_4[17];
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_4[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_12_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_12_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_5[17];
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_5[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_11_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_11_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_6[17];
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_6[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_10_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_10_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_7[17];
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_7[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_9_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_9_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_8[17];
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_8[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_8_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_8_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_9[17];
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_9[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_7_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_7_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_10[17];
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_10[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_6_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_6_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_11[17];
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_11[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_5_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_5_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_12[17];
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_12[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_4_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_4_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_13[17];
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_13[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_3_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_3_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_14[17];
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_14[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_2_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_2_sva);
      IntShiftRight_18U_2U_8U_obits_fixed_slc_data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_acc_psp_17_7_itm_3
          <= z_out_15[17];
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_IntShiftRight_18U_2U_8U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_15[0]) | IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_1_sva))
          | IntShiftRight_18U_2U_8U_obits_fixed_and_unfl_1_sva);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      o_data_data_15_6_1_sva_9 <= 6'b0;
      o_data_data_15_13_10_sva_5 <= 4'b0;
      o_data_data_15_9_7_sva_5 <= 3'b0;
      o_data_data_14_6_1_sva_9 <= 6'b0;
      o_data_data_14_13_10_sva_5 <= 4'b0;
      o_data_data_14_9_7_sva_5 <= 3'b0;
      o_data_data_13_6_1_sva_9 <= 6'b0;
      o_data_data_13_13_10_sva_5 <= 4'b0;
      o_data_data_13_9_7_sva_5 <= 3'b0;
      o_data_data_12_6_1_sva_9 <= 6'b0;
      o_data_data_12_13_10_sva_5 <= 4'b0;
      o_data_data_12_9_7_sva_5 <= 3'b0;
      o_data_data_11_6_1_sva_9 <= 6'b0;
      o_data_data_11_13_10_sva_5 <= 4'b0;
      o_data_data_11_9_7_sva_5 <= 3'b0;
      o_data_data_10_6_1_sva_9 <= 6'b0;
      o_data_data_10_13_10_sva_5 <= 4'b0;
      o_data_data_10_9_7_sva_5 <= 3'b0;
      o_data_data_9_6_1_sva_9 <= 6'b0;
      o_data_data_9_13_10_sva_5 <= 4'b0;
      o_data_data_9_9_7_sva_5 <= 3'b0;
      o_data_data_8_6_1_sva_9 <= 6'b0;
      o_data_data_8_13_10_sva_5 <= 4'b0;
      o_data_data_8_9_7_sva_5 <= 3'b0;
      o_data_data_7_6_1_sva_9 <= 6'b0;
      o_data_data_7_13_10_sva_5 <= 4'b0;
      o_data_data_7_9_7_sva_5 <= 3'b0;
      o_data_data_6_6_1_sva_9 <= 6'b0;
      o_data_data_6_13_10_sva_5 <= 4'b0;
      o_data_data_6_9_7_sva_5 <= 3'b0;
      o_data_data_5_6_1_sva_9 <= 6'b0;
      o_data_data_5_13_10_sva_5 <= 4'b0;
      o_data_data_5_9_7_sva_5 <= 3'b0;
      o_data_data_4_6_1_sva_9 <= 6'b0;
      o_data_data_4_13_10_sva_5 <= 4'b0;
      o_data_data_4_9_7_sva_5 <= 3'b0;
      o_data_data_3_6_1_sva_9 <= 6'b0;
      o_data_data_3_13_10_sva_5 <= 4'b0;
      o_data_data_3_9_7_sva_5 <= 3'b0;
      o_data_data_2_6_1_sva_9 <= 6'b0;
      o_data_data_2_13_10_sva_5 <= 4'b0;
      o_data_data_2_9_7_sva_5 <= 3'b0;
      o_data_data_1_6_1_sva_9 <= 6'b0;
      o_data_data_1_13_10_sva_5 <= 4'b0;
      o_data_data_1_9_7_sva_5 <= 3'b0;
      o_data_data_0_6_1_sva_9 <= 6'b0;
      o_data_data_0_13_10_sva_5 <= 4'b0;
      o_data_data_0_9_7_sva_5 <= 3'b0;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= 1'b0;
    end
    else if ( o_data_data_and_80_cse ) begin
      o_data_data_15_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva));
      o_data_data_15_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva));
      o_data_data_15_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva));
      o_data_data_14_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva));
      o_data_data_14_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva));
      o_data_data_14_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva));
      o_data_data_13_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva));
      o_data_data_13_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva));
      o_data_data_13_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva));
      o_data_data_12_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva));
      o_data_data_12_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva));
      o_data_data_12_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva));
      o_data_data_11_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva));
      o_data_data_11_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva));
      o_data_data_11_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva));
      o_data_data_10_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva));
      o_data_data_10_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva));
      o_data_data_10_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva));
      o_data_data_9_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva));
      o_data_data_9_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva));
      o_data_data_9_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva));
      o_data_data_8_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva));
      o_data_data_8_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva));
      o_data_data_8_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva));
      o_data_data_7_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva));
      o_data_data_7_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva));
      o_data_data_7_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva));
      o_data_data_6_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva));
      o_data_data_6_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva));
      o_data_data_6_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva));
      o_data_data_5_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva));
      o_data_data_5_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva));
      o_data_data_5_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva));
      o_data_data_4_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva));
      o_data_data_4_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva));
      o_data_data_4_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva));
      o_data_data_3_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva));
      o_data_data_3_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva));
      o_data_data_3_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva));
      o_data_data_2_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva));
      o_data_data_2_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva));
      o_data_data_2_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva));
      o_data_data_1_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva));
      o_data_data_1_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva));
      o_data_data_1_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva));
      o_data_data_0_6_1_sva_9 <= ~(MUX_v_6_2_2((data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl),
          6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva));
      o_data_data_0_13_10_sva_5 <= ~(MUX_v_4_2_2((data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl),
          4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva));
      o_data_data_0_9_7_sva_5 <= ~(MUX_v_3_2_2((data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl),
          3'b111, IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva));
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva);
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_sva);
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_15[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva);
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_15[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_15_sva);
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_14[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva);
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_14[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_14_sva);
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_13[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva);
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_13[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_13_sva);
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_12[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva);
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_12[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_12_sva);
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_11[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva);
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_11[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_11_sva);
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_10[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva);
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_10[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_10_sva);
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_9[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva);
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_9[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_9_sva);
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_8[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva);
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_8[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_8_sva);
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_7[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva);
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_7[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_7_sva);
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_6[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva);
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_6[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_6_sva);
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_5[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva);
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_5[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_5_sva);
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_4[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva);
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_4[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_4_sva);
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_3[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva);
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_3[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_3_sva);
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_2[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva);
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_2[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_2_sva);
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_itm_3
          <= ~((~((z_out_1[14]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva);
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_IntShiftRight_18U_2U_16U_obits_fixed_nor_1_itm_3
          <= ~((~((z_out_1[0]) | IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva))
          | IntShiftRight_18U_2U_16U_obits_fixed_and_unfl_1_sva);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_544_nl) ) begin
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_7 <= FpAdd_6U_10U_o_mant_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_549_nl) ) begin
      FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_7 <= FpAdd_6U_10U_1_o_mant_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_554_nl) ) begin
      FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_7 <= FpAdd_6U_10U_2_o_mant_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_559_nl) ) begin
      FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_7 <= FpAdd_6U_10U_3_o_mant_3_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_560_nl) ) begin
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_7 <= FpAdd_6U_10U_o_mant_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_563_nl) ) begin
      FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_7 <= FpAdd_6U_10U_1_o_mant_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_564_nl) ) begin
      FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_7 <= FpAdd_6U_10U_2_o_mant_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_565_nl) ) begin
      FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_7 <= FpAdd_6U_10U_3_o_mant_2_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_566_nl) ) begin
      FpAdd_6U_10U_o_mant_lpi_1_dfm_7 <= FpAdd_6U_10U_o_mant_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_567_nl) ) begin
      FpAdd_6U_10U_1_o_mant_lpi_1_dfm_7 <= FpAdd_6U_10U_1_o_mant_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_568_nl) ) begin
      FpAdd_6U_10U_2_o_mant_lpi_1_dfm_7 <= FpAdd_6U_10U_2_o_mant_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (mux_569_nl) ) begin
      FpAdd_6U_10U_3_o_mant_lpi_1_dfm_7 <= FpAdd_6U_10U_3_o_mant_lpi_1_dfm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_7 <= 10'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_2_o_mant_and_8_cse ) begin
      FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_7 <= FpAdd_6U_10U_2_o_mant_1_lpi_1_dfm_6;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_7 <= 10'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_1_o_mant_and_8_cse ) begin
      FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_7 <= FpAdd_6U_10U_1_o_mant_1_lpi_1_dfm_6;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_7 <= 10'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_o_mant_and_8_cse ) begin
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_7 <= FpAdd_6U_10U_o_mant_1_lpi_1_dfm_6;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_7 <= 10'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_3_o_mant_and_8_cse ) begin
      FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_7 <= FpAdd_6U_10U_3_o_mant_1_lpi_1_dfm_6;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_13_land_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (~ (mux_604_nl)) ) begin
      IsNaN_6U_10U_13_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_13_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (~ (mux_605_nl)) ) begin
      IsNaN_6U_10U_13_land_1_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_13_land_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_64) & (~ (mux_606_nl)) ) begin
      IsNaN_6U_10U_13_land_lpi_1_dfm_4 <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1348_rgt | and_1351_rgt | and_1354_rgt | and_1357_rgt)
        & mux_11_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[185:176]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          (chn_data_in_rsci_d_mxwt[57:48]), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_6_mx0w4,
          {and_1348_rgt , and_1351_rgt , and_1354_rgt , and_1357_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_5 <= MUX_v_2_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3, and_dcpl_1074);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w2, and_dcpl_1074);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm <= IsNaN_6U_10U_1_IsNaN_6U_10U_1_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1362_rgt | and_1365_rgt | and_1368_rgt | and_1371_rgt)
        & mux_24_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[121:112]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          (chn_data_in_rsci_d_mxwt[185:176]), FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          {and_1362_rgt , and_1365_rgt , and_1368_rgt , and_1371_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_25_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_1075) | and_1373_rgt) & mux_24_cse
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0, and_1373_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm <= IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1376_rgt | and_1379_rgt | and_1382_rgt | and_1385_rgt)
        & mux_33_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[185:176]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_4_FpExpoWidthInc_5U_6U_10U_1U_1U_4_or_6_mx0w1,
          (chn_data_in_rsci_d_mxwt[121:112]), FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          {and_1376_rgt , and_1379_rgt , and_1382_rgt , and_1385_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_6 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_and_21_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0, and_dcpl_1102);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_1_1 <= MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]), and_dcpl_1102);
      FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_expo_5_4_lpi_1_dfm_3_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          and_dcpl_1102);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm <= IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & (and_1390_rgt | and_1393_rgt | and_1396_rgt | and_1399_rgt)
        & mux_46_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_4_2((chn_data_in_rsci_d_mxwt[121:112]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_6_FpExpoWidthInc_5U_6U_10U_1U_1U_6_or_6_mx0w1,
          (chn_data_in_rsci_d_mxwt[249:240]), FpExpoWidthInc_5U_6U_10U_1U_1U_7_FpExpoWidthInc_5U_6U_10U_1U_1U_7_or_6_mx0w4,
          {and_1390_rgt , and_1393_rgt , and_1396_rgt , and_1399_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_6 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_74 & and_dcpl_1103) | and_1401_rgt) & mux_46_cse
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_6 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_3_0_lpi_1_dfm_3_mx0w2, and_1401_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & (~ or_dcpl_303) & (mux_48_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_5 <= FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_23 | or_dcpl_21 | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp
        | (fsm_output[0]))) ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm <= IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_0_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_and_22_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1];
      FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_expo_5_4_lpi_1_dfm_3_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_610_nl) ) begin
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_4,
          FpAdd_6U_10U_4_mux_45_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_612_nl) ) begin
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_4,
          FpAdd_6U_10U_4_mux_13_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_613_nl) ) begin
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_4,
          FpAdd_6U_10U_5_mux_45_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_615_nl) ) begin
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_4,
          FpAdd_6U_10U_5_mux_13_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_616_nl) ) begin
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_4,
          FpAdd_6U_10U_6_mux_45_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_618_nl) ) begin
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_4,
          FpAdd_6U_10U_6_mux_13_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_619_nl) ) begin
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_4,
          FpAdd_6U_10U_4_mux_29_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_620_nl) ) begin
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_4,
          FpAdd_6U_10U_5_mux_29_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_621_nl) ) begin
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_4,
          FpAdd_6U_10U_6_mux_29_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_624_nl) ) begin
      FpAdd_6U_10U_1_o_sign_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_sign_lpi_1_dfm_4,
          FpAdd_6U_10U_4_mux_61_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_626_nl) ) begin
      FpAdd_6U_10U_2_o_sign_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_2_o_sign_lpi_1_dfm_4,
          FpAdd_6U_10U_5_mux_61_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_628_nl) ) begin
      FpAdd_6U_10U_3_o_sign_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_3_o_sign_lpi_1_dfm_4,
          FpAdd_6U_10U_6_mux_61_mx1w1, and_dcpl_1122);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_nor_1_itm_2 <= 1'b0;
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_cse ) begin
      IsNaN_6U_10U_9_nor_1_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_nor_1_tmp, IsNaN_6U_10U_9_nor_1_itm,
          and_dcpl_78);
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp,
          IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_nor_2_itm_2 <= 1'b0;
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_7_cse ) begin
      IsNaN_6U_10U_9_nor_2_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_nor_2_tmp, IsNaN_6U_10U_9_nor_2_itm,
          and_dcpl_78);
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp,
          IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_nor_3_itm_2 <= 1'b0;
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_9_cse ) begin
      IsNaN_6U_10U_9_nor_3_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_nor_3_tmp, IsNaN_6U_10U_9_nor_3_itm,
          and_dcpl_78);
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp,
          IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_13_nor_1_itm_2 <= 1'b0;
      IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_13_and_cse ) begin
      IsNaN_6U_10U_13_nor_1_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_10_nor_1_tmp, IsNaN_6U_10U_13_nor_1_itm,
          and_dcpl_78);
      IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2 <= MUX_s_1_2_2(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp,
          IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm, and_dcpl_78);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_18U_2U_16U_mbits_fixed_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_1_20_2_1 <= 19'b0;
    end
    else if ( IntShiftRight_18U_2U_16U_mbits_fixed_and_cse ) begin
      IntShiftRight_18U_2U_16U_mbits_fixed_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_15_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_14_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_13_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_12_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_11_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_10_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_9_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_8_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_7_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_6_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_5_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_4_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_3_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_2_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_16U_mbits_fixed_1_tmp, IntShiftRight_18U_2U_16U_mbits_fixed_and_31_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_18U_2U_16U_obits_fixed_and_80_cse ) begin
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm, and_dcpl_1126);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_18U_2U_8U_mbits_fixed_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_15_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_14_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_13_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_12_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_11_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_10_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_9_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_8_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_7_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_6_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_5_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_4_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_3_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_2_sva_1_20_2_1 <= 19'b0;
      IntShiftRight_18U_2U_8U_mbits_fixed_1_sva_1_20_2_1 <= 19'b0;
    end
    else if ( IntShiftRight_18U_2U_8U_mbits_fixed_and_cse ) begin
      IntShiftRight_18U_2U_8U_mbits_fixed_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_15_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_15_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_14_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_14_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_13_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_13_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_12_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_12_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_11_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_11_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_10_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_10_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_9_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_9_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_8_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_8_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_7_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_7_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_6_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_6_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_5_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_5_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_4_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_4_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_3_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_3_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_2_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_2_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
      IntShiftRight_18U_2U_8U_mbits_fixed_1_sva_1_20_2_1 <= MUX_v_19_2_2((IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[20:2]),
          reg_IntShiftRight_18U_2U_8U_mbits_fixed_1_tmp, IntShiftRight_18U_2U_8U_mbits_fixed_and_31_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( IntShiftRight_18U_2U_8U_obits_fixed_and_144_cse ) begin
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2 <= MUX_s_1_2_2(data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0,
          data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm, and_dcpl_1129);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_640_nl) ) begin
      FpAdd_6U_10U_7_o_sign_1_lpi_1_dfm_2 <= MUX_s_1_2_2(FpAdd_6U_10U_7_mux_13_mx1w0,
          FpAdd_6U_10U_o_sign_1_lpi_1_dfm_4, and_dcpl_1119);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_641_nl) ) begin
      FpAdd_6U_10U_7_o_sign_2_lpi_1_dfm_2 <= MUX_s_1_2_2(FpAdd_6U_10U_7_mux_29_mx1w0,
          FpAdd_6U_10U_o_sign_2_lpi_1_dfm_4, and_dcpl_1119);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_642_nl) ) begin
      FpAdd_6U_10U_7_o_sign_3_lpi_1_dfm_2 <= MUX_s_1_2_2(FpAdd_6U_10U_7_mux_45_mx1w0,
          FpAdd_6U_10U_o_sign_3_lpi_1_dfm_4, and_dcpl_1119);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_3_b_int_mant_p1_and_cse & FpAdd_6U_10U_1_o_sign_FpAdd_6U_10U_1_o_sign_or_7_cse
        & (mux_644_nl) ) begin
      FpAdd_6U_10U_7_o_sign_lpi_1_dfm_2 <= MUX_s_1_2_2(FpAdd_6U_10U_7_mux_61_mx1w0,
          FpAdd_6U_10U_o_sign_lpi_1_dfm_4, and_dcpl_1119);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_sign_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_IsNaN_6U_10U_and_tmp) | (FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_tmp
        & FpAdd_6U_10U_o_sign_1_lpi_1_dfm_3_mx0c2) | FpAdd_6U_10U_o_sign_or_1_rgt)
        & mux_tmp_49 ) begin
      FpAdd_6U_10U_o_sign_1_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[15]),
          (~ (chn_data_in_rsci_d_mxwt[143])), FpAdd_6U_10U_o_sign_or_1_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp) |
        (FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_tmp & FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_3_mx0c2)
        | FpAdd_6U_10U_1_o_sign_or_1_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_1_o_sign_1_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[79]),
          (chn_data_in_rsci_d_mxwt[143]), FpAdd_6U_10U_1_o_sign_or_1_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm <= 1'b0;
      IsNaN_6U_10U_9_nor_1_itm <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_11_cse ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_itm <= IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp;
      IsNaN_6U_10U_9_nor_1_itm <= IsNaN_6U_10U_9_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_tmp) |
        (FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_tmp & FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_3_mx0c2)
        | m_row1_if_d2_or_1_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_2_o_sign_1_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[143]),
          (~ (chn_data_in_rsci_d_mxwt[79])), m_row1_if_d2_or_1_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm <= 1'b0;
      IsNaN_6U_10U_9_nor_2_itm <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_13_cse ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_itm <= IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp;
      IsNaN_6U_10U_9_nor_2_itm <= IsNaN_6U_10U_9_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp) |
        (FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_tmp & FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_3_mx0c2)
        | FpAdd_6U_10U_1_o_sign_or_4_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_3_o_sign_1_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[79]),
          (~ (chn_data_in_rsci_d_mxwt[207])), FpAdd_6U_10U_1_o_sign_or_4_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm <= 1'b0;
      IsNaN_6U_10U_9_nor_3_itm <= 1'b0;
    end
    else if ( IsNaN_6U_10U_9_and_15_cse ) begin
      IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_itm <= IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp;
      IsNaN_6U_10U_9_nor_3_itm <= IsNaN_6U_10U_9_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_sign_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_IsNaN_6U_10U_and_1_tmp) | (FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_1_tmp
        & and_1439_m1c) | FpAdd_6U_10U_o_sign_or_11_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_o_sign_2_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[31]),
          (~ (chn_data_in_rsci_d_mxwt[159])), FpAdd_6U_10U_o_sign_or_11_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (and_1440_rgt | and_1442_rgt | and_1444_rgt) & mux_tmp_49
        ) begin
      FpAdd_6U_10U_1_o_sign_2_lpi_1_dfm_4 <= MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[95]),
          (chn_data_in_rsci_d_mxwt[159]), FpAdd_6U_10U_1_mux_19_mx0w2, {and_1440_rgt
          , and_1442_rgt , and_1444_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_1_tmp)
        | (FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_1_tmp & and_1449_m1c)
        | m_row1_if_d2_or_11_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_2_o_sign_2_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[159]),
          (~ (chn_data_in_rsci_d_mxwt[95])), m_row1_if_d2_or_11_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp)
        | (FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_1_tmp & and_1454_m1c)
        | FpAdd_6U_10U_1_o_sign_or_17_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_3_o_sign_2_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[95]),
          (~ (chn_data_in_rsci_d_mxwt[223])), FpAdd_6U_10U_1_o_sign_or_17_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_sign_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_IsNaN_6U_10U_and_2_tmp) | (FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_2_tmp
        & and_1459_m1c) | FpAdd_6U_10U_o_sign_or_8_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_o_sign_3_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[47]),
          (~ (chn_data_in_rsci_d_mxwt[175])), FpAdd_6U_10U_o_sign_or_8_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (and_1460_rgt | and_1462_rgt | and_1464_rgt) & mux_tmp_49
        ) begin
      FpAdd_6U_10U_1_o_sign_3_lpi_1_dfm_4 <= MUX1HOT_s_1_3_2((chn_data_in_rsci_d_mxwt[111]),
          (chn_data_in_rsci_d_mxwt[175]), FpAdd_6U_10U_1_mux_36_mx0w2, {and_1460_rgt
          , and_1462_rgt , and_1464_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm <= 1'b0;
      IsNaN_6U_10U_13_nor_1_itm <= 1'b0;
    end
    else if ( IsNaN_6U_10U_13_and_3_cse ) begin
      IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm <= IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp;
      IsNaN_6U_10U_13_nor_1_itm <= IsNaN_6U_10U_10_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_2_tmp)
        | (FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_2_tmp & and_1469_m1c)
        | m_row1_if_d2_or_8_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_2_o_sign_3_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[175]),
          (~ (chn_data_in_rsci_d_mxwt[111])), m_row1_if_d2_or_8_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp)
        | (FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_2_tmp & and_1474_m1c)
        | FpAdd_6U_10U_1_o_sign_or_14_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_3_o_sign_3_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[111]),
          (~ (chn_data_in_rsci_d_mxwt[239])), FpAdd_6U_10U_1_o_sign_or_14_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_3_o_sign_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp)
        | (FpAdd_6U_10U_3_is_a_greater_FpAdd_6U_10U_3_is_a_greater_or_3_tmp & FpAdd_6U_10U_3_o_sign_lpi_1_dfm_3_mx0c2)
        | FpAdd_6U_10U_1_o_sign_or_9_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_3_o_sign_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[127]),
          (~ (chn_data_in_rsci_d_mxwt[255])), FpAdd_6U_10U_1_o_sign_or_9_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_2_o_sign_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_4_IsNaN_6U_10U_4_and_3_tmp)
        | (FpAdd_6U_10U_2_is_a_greater_FpAdd_6U_10U_2_is_a_greater_or_3_tmp & FpAdd_6U_10U_2_o_sign_lpi_1_dfm_3_mx0c2)
        | m_row1_if_d2_or_3_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_2_o_sign_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[191]),
          (~ (chn_data_in_rsci_d_mxwt[127])), m_row1_if_d2_or_3_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_sign_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp)
        | (FpAdd_6U_10U_1_is_a_greater_FpAdd_6U_10U_1_is_a_greater_or_3_tmp & FpAdd_6U_10U_1_o_sign_lpi_1_dfm_3_mx0c2)
        | FpAdd_6U_10U_1_o_sign_or_6_rgt) & mux_tmp_49 ) begin
      FpAdd_6U_10U_1_o_sign_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[127]),
          (chn_data_in_rsci_d_mxwt[191]), FpAdd_6U_10U_1_o_sign_or_6_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_sign_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_181_cse & IsNaN_6U_10U_IsNaN_6U_10U_and_3_tmp) | (FpAdd_6U_10U_is_a_greater_FpAdd_6U_10U_is_a_greater_or_3_tmp
        & FpAdd_6U_10U_o_sign_lpi_1_dfm_3_mx0c2) | FpAdd_6U_10U_o_sign_or_3_rgt)
        & mux_tmp_49 ) begin
      FpAdd_6U_10U_o_sign_lpi_1_dfm_4 <= MUX_s_1_2_2((chn_data_in_rsci_d_mxwt[63]),
          (~ (chn_data_in_rsci_d_mxwt[191])), FpAdd_6U_10U_o_sign_or_3_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= 1'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_1_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_2_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_3_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_4_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_5_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_6_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_7_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_8_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_9_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_10_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_11_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_12_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_13_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_14_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_15_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_tmp <= 19'b0;
    end
    else if ( IntShiftRight_18U_2U_16U_obits_fixed_and_cse ) begin
      data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm <= data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_1_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_2_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_3_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_4_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_5_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_6_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_7_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_8_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_9_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_10_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_11_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_12_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_13_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_14_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_15_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_16U_mbits_fixed_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[20:2];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= 1'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_1_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_2_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_3_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_4_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_5_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_6_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_7_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_8_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_9_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_10_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_11_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_12_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_13_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_14_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_15_tmp <= 19'b0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_tmp <= 19'b0;
    end
    else if ( IntShiftRight_18U_2U_8U_obits_fixed_and_cse ) begin
      data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm <= data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_mx0w0;
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_1_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_2_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_3_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_4_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_5_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_6_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_7_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_8_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_9_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_10_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_11_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_12_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_13_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_14_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_15_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_mx0w0[20:2];
      reg_IntShiftRight_18U_2U_8U_mbits_fixed_tmp <= IntShiftRight_18U_2U_16U_mbits_fixed_sva_mx0w0[20:2];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSubExt_16U_16U_17U_2_o_acc_2_itm <= 17'b0;
      IntSubExt_16U_16U_17U_1_o_acc_2_itm <= 17'b0;
      IntAddExt_16U_16U_17U_o_acc_1_itm <= 17'b0;
      IntSubExt_16U_16U_17U_o_acc_2_itm <= 17'b0;
      IntSubExt_16U_16U_17U_2_o_acc_1_itm <= 17'b0;
      IntSubExt_16U_16U_17U_1_o_acc_1_itm <= 17'b0;
      IntAddExt_16U_16U_17U_o_acc_itm <= 17'b0;
      IntSubExt_16U_16U_17U_o_acc_1_itm <= 17'b0;
      m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva <= 17'b0;
      m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva <= 17'b0;
      m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva <= 17'b0;
      m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva <= 17'b0;
      m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva <= 17'b0;
      m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva <= 17'b0;
      m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva <= 17'b0;
      m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva <= 17'b0;
    end
    else if ( IntSubExt_16U_16U_17U_2_o_and_cse ) begin
      IntSubExt_16U_16U_17U_2_o_acc_2_itm <= IntSubExt_16U_16U_17U_2_o_acc_2_itm_mx0w0;
      IntSubExt_16U_16U_17U_1_o_acc_2_itm <= IntSubExt_16U_16U_17U_1_o_acc_2_itm_mx0w0;
      IntAddExt_16U_16U_17U_o_acc_1_itm <= IntAddExt_16U_16U_17U_o_acc_1_itm_mx0w0;
      IntSubExt_16U_16U_17U_o_acc_2_itm <= IntSubExt_16U_16U_17U_o_acc_2_itm_mx0w0;
      IntSubExt_16U_16U_17U_2_o_acc_1_itm <= IntSubExt_16U_16U_17U_2_o_acc_1_itm_mx0w0;
      IntSubExt_16U_16U_17U_1_o_acc_1_itm <= IntSubExt_16U_16U_17U_1_o_acc_1_itm_mx0w0;
      IntAddExt_16U_16U_17U_o_acc_itm <= IntAddExt_16U_16U_17U_o_acc_itm_mx0w0;
      IntSubExt_16U_16U_17U_o_acc_1_itm <= IntSubExt_16U_16U_17U_o_acc_1_itm_mx0w0;
      m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva <= m_row3_3_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
      m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva <= m_row3_2_IntSubExt_16U_16U_17U_2_o_acc_ncse_sva_mx0w0;
      m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva <= m_row2_3_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
      m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva <= m_row2_2_IntSubExt_16U_16U_17U_1_o_acc_ncse_sva_mx0w0;
      m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva <= m_row1_3_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
      m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva <= m_row1_2_IntAddExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
      m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva <= m_row0_3_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
      m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva <= m_row0_2_IntSubExt_16U_16U_17U_o_acc_ncse_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_cse ) begin
      reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4[1]), FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_1,
          {and_dcpl_823 , and_dcpl_824 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_lpi_1_dfm_4[0]), FpAdd_6U_10U_3_qr_5_4_lpi_1_dfm_0,
          {and_dcpl_823 , and_dcpl_824 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4[1]), FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_1,
          {and_dcpl_833 , and_dcpl_834 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_3_lpi_1_dfm_4[0]), FpAdd_6U_10U_3_qr_5_4_3_lpi_1_dfm_0,
          {and_dcpl_833 , and_dcpl_834 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4[1]), FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_1,
          {and_dcpl_843 , and_dcpl_844 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_2_lpi_1_dfm_4[0]), FpAdd_6U_10U_3_qr_5_4_2_lpi_1_dfm_0,
          {and_dcpl_843 , and_dcpl_844 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4[1]), FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_1,
          {and_dcpl_853 , and_dcpl_854 , or_dcpl_1});
      reg_FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          (FpExpoWidthInc_5U_6U_10U_1U_1U_7_o_expo_5_4_1_lpi_1_dfm_4[0]), FpAdd_6U_10U_3_qr_5_4_1_lpi_1_dfm_0,
          {and_dcpl_853 , and_dcpl_854 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]), FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_1,
          {and_dcpl_863 , and_dcpl_864 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_6_psp,
          FpAdd_6U_10U_2_qr_5_4_lpi_1_dfm_0, {and_dcpl_863 , and_dcpl_864 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]), FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_1,
          {and_dcpl_873 , and_dcpl_874 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_4_psp,
          FpAdd_6U_10U_2_qr_5_4_3_lpi_1_dfm_0, {and_dcpl_873 , and_dcpl_874 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]), FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_1,
          {and_dcpl_883 , and_dcpl_884 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_2_psp,
          FpAdd_6U_10U_2_qr_5_4_2_lpi_1_dfm_0, {and_dcpl_883 , and_dcpl_884 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]), FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_1,
          {and_dcpl_893 , and_dcpl_894 , or_dcpl_1});
      reg_FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_5_if_3_or_psp,
          FpAdd_6U_10U_2_qr_5_4_1_lpi_1_dfm_0, {and_dcpl_893 , and_dcpl_894 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]), FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_1,
          {and_dcpl_903 , and_dcpl_904 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_6_psp,
          FpAdd_6U_10U_1_qr_5_4_lpi_1_dfm_0, {and_dcpl_903 , and_dcpl_904 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]), FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_1,
          {and_dcpl_913 , and_dcpl_914 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_4_psp,
          FpAdd_6U_10U_1_qr_5_4_3_lpi_1_dfm_0, {and_dcpl_913 , and_dcpl_914 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]), FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_1,
          {and_dcpl_923 , and_dcpl_924 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_2_psp,
          FpAdd_6U_10U_1_qr_5_4_2_lpi_1_dfm_0, {and_dcpl_923 , and_dcpl_924 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]), FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_1,
          {and_dcpl_933 , and_dcpl_934 , or_dcpl_1});
      reg_FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_4[0]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_3_or_psp,
          FpAdd_6U_10U_1_qr_5_4_1_lpi_1_dfm_0, {and_dcpl_933 , and_dcpl_934 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[1]), FpAdd_6U_10U_qr_5_4_lpi_1_dfm_1,
          {and_dcpl_943 , and_dcpl_944 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_4[0]), FpAdd_6U_10U_qr_5_4_lpi_1_dfm_0,
          {and_dcpl_943 , and_dcpl_944 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[1]), FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_1,
          {and_dcpl_953 , and_dcpl_954 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_4[0]), FpAdd_6U_10U_qr_5_4_3_lpi_1_dfm_0,
          {and_dcpl_953 , and_dcpl_954 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[1]), FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_1,
          {and_dcpl_963 , and_dcpl_964 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_4[0]), FpAdd_6U_10U_qr_5_4_2_lpi_1_dfm_0,
          {and_dcpl_963 , and_dcpl_964 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3[1]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[1]), FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_1,
          {and_dcpl_973 , and_dcpl_974 , or_dcpl_1});
      reg_FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3[0]),
          (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_4[0]), FpAdd_6U_10U_qr_5_4_1_lpi_1_dfm_0,
          {and_dcpl_973 , and_dcpl_974 , or_dcpl_1});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_3_o_expo_and_13_ssc ) begin
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_3_o_expo_and_12_ssc ) begin
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_3_o_expo_and_11_ssc ) begin
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_o_expo_and_13_ssc ) begin
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_1_o_expo_and_13_ssc ) begin
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_2_o_expo_and_13_ssc ) begin
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_o_expo_and_12_ssc ) begin
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_1_o_expo_and_12_ssc ) begin
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_2_o_expo_and_12_ssc ) begin
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_o_expo_and_11_ssc ) begin
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_1_o_expo_and_11_ssc ) begin
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_2_o_expo_and_11_ssc ) begin
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp <= reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_1 <= reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1;
      reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_10_tmp_2 <= reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_38_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp, FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_6_qr_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_38_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_5_qr_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_38_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_4_qr_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_42_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp,
          {and_777_rgt , and_779_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_1,
          {and_777_rgt , and_779_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_6_qr_lpi_1_dfm_tmp_2,
          {and_777_rgt , and_779_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_42_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp,
          {and_761_rgt , and_763_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_1,
          {and_761_rgt , and_763_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_5_qr_lpi_1_dfm_tmp_2,
          {and_761_rgt , and_763_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_42_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp,
          {and_745_rgt , and_747_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_1,
          {and_745_rgt , and_747_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_3_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_4_qr_lpi_1_dfm_tmp_2,
          {and_745_rgt , and_747_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_38_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp, FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_7_qr_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_42_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp,
          {and_793_rgt , and_795_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_1,
          {and_793_rgt , and_795_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_3_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_3_o_expo_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_7_qr_lpi_1_dfm_tmp_2,
          {and_793_rgt , and_795_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_35_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp, FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_6_qr_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_35_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_5_qr_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_35_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_4_qr_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_39_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp,
          {and_765_rgt , and_767_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_1,
          {and_765_rgt , and_767_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_6_qr_2_lpi_1_dfm_tmp_2,
          {and_765_rgt , and_767_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_39_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp,
          {and_749_rgt , and_751_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_1,
          {and_749_rgt , and_751_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_5_qr_2_lpi_1_dfm_tmp_2,
          {and_749_rgt , and_751_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_39_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp,
          {and_733_rgt , and_735_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_1,
          {and_733_rgt , and_735_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_4_qr_2_lpi_1_dfm_tmp_2,
          {and_733_rgt , and_735_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_36_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp, FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_6_qr_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_36_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_5_qr_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_36_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_4_qr_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_40_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp,
          {and_769_rgt , and_771_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_1,
          {and_769_rgt , and_771_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_6_qr_3_lpi_1_dfm_tmp_2,
          {and_769_rgt , and_771_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_40_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp,
          {and_753_rgt , and_755_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_1,
          {and_753_rgt , and_755_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_5_qr_3_lpi_1_dfm_tmp_2,
          {and_753_rgt , and_755_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_40_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp,
          {and_737_rgt , and_739_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_1,
          {and_737_rgt , and_739_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_4_qr_3_lpi_1_dfm_tmp_2,
          {and_737_rgt , and_739_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_37_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp, FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_6_qr_4_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_37_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_5_qr_4_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_37_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp, FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_4_qr_4_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_6_and_41_ssc ) begin
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp,
          {and_773_rgt , and_775_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_1,
          {and_773_rgt , and_775_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_6_qr_4_lpi_1_dfm_tmp_2,
          {and_773_rgt , and_775_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_5_and_41_ssc ) begin
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp,
          {and_757_rgt , and_759_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_1,
          {and_757_rgt , and_759_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_5_qr_4_lpi_1_dfm_tmp_2,
          {and_757_rgt , and_759_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_4_and_41_ssc ) begin
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp,
          {and_741_rgt , and_743_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_1,
          {and_741_rgt , and_743_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_2_o_expo_1_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_3_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_4_qr_4_lpi_1_dfm_tmp_2,
          {and_741_rgt , and_743_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_35_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp, FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_7_qr_2_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_39_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp,
          {and_781_rgt , and_783_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_1,
          {and_781_rgt , and_783_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_o_expo_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_7_qr_2_lpi_1_dfm_tmp_2,
          {and_781_rgt , and_783_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_36_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp, FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_7_qr_3_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_40_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp,
          {and_785_rgt , and_787_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_1,
          {and_785_rgt , and_787_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_1_o_expo_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_7_qr_3_lpi_1_dfm_tmp_2,
          {and_785_rgt , and_787_rgt , and_dcpl_78});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_37_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp, FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_1 <= MUX_s_1_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1, FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1);
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_2 <= MUX_v_4_2_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2, FpAdd_6U_10U_7_qr_4_lpi_1_dfm_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1 <= 1'b0;
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2 <= 4'b0;
    end
    else if ( FpAdd_6U_10U_7_and_41_ssc ) begin
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp, reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp,
          {and_789_rgt , and_791_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_1,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_1, reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_1,
          {and_789_rgt , and_791_rgt , and_dcpl_78});
      reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_2_tmp_2 <= MUX1HOT_v_4_3_2(reg_FpAdd_6U_10U_2_o_expo_2_lpi_1_dfm_9_tmp_2,
          reg_FpAdd_6U_10U_2_o_expo_lpi_1_dfm_9_tmp_2, reg_FpAdd_6U_10U_7_qr_4_lpi_1_dfm_tmp_2,
          {and_789_rgt , and_791_rgt , and_dcpl_78});
    end
  end
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_6_nl = MUX_v_4_2_2(({3'b0 ,
      (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_1_sva[10])}), (FpAdd_6U_10U_4_o_expo_1_lpi_2[3:0]),
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_255_nl = ~ data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_2_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_6_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_255_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_172_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_2_nl),
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_1_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_172_nl), 4'b1111, IsNaN_6U_10U_16_land_1_lpi_1_dfm_3);
  assign or_1299_nl = or_dcpl_203 | data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_1_nl = MUX_s_1_2_2(data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1299_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_1_nl = MUX_s_1_2_2(data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_203);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_nl
      = ((~ (FpAdd_6U_10U_4_o_expo_1_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_1_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_1_nl))) | (~ data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_1_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_17_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_2_sva[10])}), (FpAdd_6U_10U_5_o_expo_1_lpi_2[3:0]),
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_256_nl = ~ data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_5_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_17_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_256_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_17_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_5_nl),
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_3_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_17_nl), 4'b1111, IsNaN_6U_10U_16_land_2_lpi_1_dfm_3);
  assign or_1305_nl = or_dcpl_209 | data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_3_nl = MUX_s_1_2_2(data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1305_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_3_nl = MUX_s_1_2_2(data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_209);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_2_nl
      = ((~ (FpAdd_6U_10U_5_o_expo_1_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_3_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_3_nl))) | (~ data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_2_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_28_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_3_sva[10])}), (FpAdd_6U_10U_6_o_expo_1_lpi_2[3:0]),
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_257_nl = ~ data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_8_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_28_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_257_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_28_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_8_nl),
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_5_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_28_nl), 4'b1111, IsNaN_6U_10U_16_land_3_lpi_1_dfm_3);
  assign or_1311_nl = or_dcpl_215 | data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_5_nl = MUX_s_1_2_2(data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1311_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_5_nl = MUX_s_1_2_2(data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_215);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_4_nl
      = ((~ (FpAdd_6U_10U_6_o_expo_1_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_5_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_5_nl))) | (~ data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_3_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_39_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_4_sva[10])}), (FpAdd_6U_10U_7_o_expo_1_lpi_2[3:0]),
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_258_nl = ~ data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_11_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_39_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_258_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_39_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_11_nl),
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_7_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_39_nl), 4'b1111, IsNaN_6U_10U_16_land_4_lpi_1_dfm_3);
  assign or_1317_nl = or_dcpl_221 | data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_7_nl = MUX_s_1_2_2(data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1317_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_7_nl = MUX_s_1_2_2(data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_221);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_6_nl
      = ((~ (FpAdd_6U_10U_7_o_expo_1_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_7_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_7_nl))) | (~ data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_4_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_50_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_5_sva[10])}), (FpAdd_6U_10U_4_o_expo_2_lpi_2[3:0]),
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_259_nl = ~ data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_14_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_50_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_259_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_50_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_14_nl),
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_9_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_50_nl), 4'b1111, IsNaN_6U_10U_16_land_5_lpi_1_dfm_3);
  assign or_1323_nl = or_dcpl_227 | data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_9_nl = MUX_s_1_2_2(data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1323_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_9_nl = MUX_s_1_2_2(data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_227);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_8_nl
      = ((~ (FpAdd_6U_10U_4_o_expo_2_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_9_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_9_nl))) | (~ data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_5_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_61_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_6_sva[10])}), (FpAdd_6U_10U_5_o_expo_2_lpi_2[3:0]),
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_260_nl = ~ data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_17_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_61_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_260_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_61_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_17_nl),
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_11_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_61_nl), 4'b1111, IsNaN_6U_10U_16_land_6_lpi_1_dfm_3);
  assign or_1329_nl = or_dcpl_233 | data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_11_nl = MUX_s_1_2_2(data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1329_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_11_nl = MUX_s_1_2_2(data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_233);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_10_nl
      = ((~ (FpAdd_6U_10U_5_o_expo_2_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_11_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_11_nl))) | (~ data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_6_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_72_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_7_sva[10])}), (FpAdd_6U_10U_6_o_expo_2_lpi_2[3:0]),
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_261_nl = ~ data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_20_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_72_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_261_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_72_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_20_nl),
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_13_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_72_nl), 4'b1111, IsNaN_6U_10U_16_land_7_lpi_1_dfm_3);
  assign or_1335_nl = or_dcpl_239 | data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_13_nl = MUX_s_1_2_2(data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1335_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_13_nl = MUX_s_1_2_2(data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_239);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_12_nl
      = ((~ (FpAdd_6U_10U_6_o_expo_2_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_13_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_13_nl))) | (~ data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_7_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_83_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_8_sva[10])}), (FpAdd_6U_10U_7_o_expo_2_lpi_2[3:0]),
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_262_nl = ~ data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_23_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_83_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_262_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_83_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_23_nl),
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_15_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_83_nl), 4'b1111, IsNaN_6U_10U_16_land_8_lpi_1_dfm_3);
  assign or_1341_nl = or_dcpl_245 | data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_15_nl = MUX_s_1_2_2(data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1341_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_15_nl = MUX_s_1_2_2(data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_245);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_14_nl
      = ((~ (FpAdd_6U_10U_7_o_expo_2_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_15_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_15_nl))) | (~ data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_8_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_94_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_9_sva[10])}), (FpAdd_6U_10U_4_o_expo_3_lpi_2[3:0]),
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_263_nl = ~ data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_26_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_94_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_263_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_94_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_26_nl),
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_17_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_94_nl), 4'b1111, IsNaN_6U_10U_16_land_9_lpi_1_dfm_3);
  assign or_1347_nl = or_dcpl_251 | data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_17_nl = MUX_s_1_2_2(data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1347_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_17_nl = MUX_s_1_2_2(data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_251);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_16_nl
      = ((~ (FpAdd_6U_10U_4_o_expo_3_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_17_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_17_nl))) | (~ data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_9_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_105_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_10_sva[10])}), (FpAdd_6U_10U_5_o_expo_3_lpi_2[3:0]),
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_264_nl = ~ data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_29_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_105_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_264_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_105_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_29_nl),
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_19_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_105_nl), 4'b1111, IsNaN_6U_10U_16_land_10_lpi_1_dfm_3);
  assign or_1353_nl = or_dcpl_257 | data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_19_nl = MUX_s_1_2_2(data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1353_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_19_nl = MUX_s_1_2_2(data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_257);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_18_nl
      = ((~ (FpAdd_6U_10U_5_o_expo_3_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_19_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_19_nl))) | (~ data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_10_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_116_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_11_sva[10])}), (FpAdd_6U_10U_6_o_expo_3_lpi_2[3:0]),
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_265_nl = ~ data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_32_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_116_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_265_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_116_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_32_nl),
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_21_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_116_nl), 4'b1111, IsNaN_6U_10U_16_land_11_lpi_1_dfm_3);
  assign or_1359_nl = or_dcpl_263 | data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_21_nl = MUX_s_1_2_2(data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1359_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_21_nl = MUX_s_1_2_2(data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_263);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_20_nl
      = ((~ (FpAdd_6U_10U_6_o_expo_3_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_21_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_21_nl))) | (~ data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_11_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_127_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_12_sva[10])}), (FpAdd_6U_10U_7_o_expo_3_lpi_2[3:0]),
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_266_nl = ~ data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_35_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_127_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_266_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_127_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_35_nl),
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_23_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_127_nl), 4'b1111, IsNaN_6U_10U_16_land_12_lpi_1_dfm_3);
  assign or_1365_nl = or_dcpl_269 | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_23_nl = MUX_s_1_2_2(data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1365_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_23_nl = MUX_s_1_2_2(data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_269);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_22_nl
      = ((~ (FpAdd_6U_10U_7_o_expo_3_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_23_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_23_nl))) | (~ data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_12_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_138_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_13_sva[10])}), (FpAdd_6U_10U_4_o_expo_lpi_2[3:0]),
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_267_nl = ~ data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_38_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_138_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_267_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_138_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_38_nl),
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_25_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_138_nl), 4'b1111, IsNaN_6U_10U_16_land_13_lpi_1_dfm);
  assign or_1371_nl = or_dcpl_275 | data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_25_nl = MUX_s_1_2_2(data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1371_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_25_nl = MUX_s_1_2_2(data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_275);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_24_nl
      = ((~ (FpAdd_6U_10U_4_o_expo_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_25_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_25_nl))) | (~ data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_13_lpi_1_dfm;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_149_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_14_sva[10])}), (FpAdd_6U_10U_5_o_expo_lpi_2[3:0]),
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_268_nl = ~ data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_41_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_149_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_268_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_149_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_41_nl),
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_27_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_149_nl), 4'b1111, IsNaN_6U_10U_16_land_14_lpi_1_dfm_3);
  assign or_1377_nl = or_dcpl_281 | data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_27_nl = MUX_s_1_2_2(data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1377_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_27_nl = MUX_s_1_2_2(data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_281);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_26_nl
      = ((~ (FpAdd_6U_10U_5_o_expo_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_27_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_27_nl))) | (~ data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_14_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_160_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_15_sva[10])}), (FpAdd_6U_10U_6_o_expo_lpi_2[3:0]),
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_269_nl = ~ data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_44_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_160_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_269_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_160_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_44_nl),
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_29_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_160_nl), 4'b1111, IsNaN_6U_10U_16_land_15_lpi_1_dfm_3);
  assign or_1383_nl = or_dcpl_287 | data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_29_nl = MUX_s_1_2_2(data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1383_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_29_nl = MUX_s_1_2_2(data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_287);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_28_nl
      = ((~ (FpAdd_6U_10U_6_o_expo_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_29_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_29_nl))) | (~ data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_15_lpi_1_dfm_3;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_171_nl = MUX_v_4_2_2(({3'b0
      , (FpMantDecShiftRight_10U_6U_10U_o_mant_sum_sva[10])}), (FpAdd_6U_10U_7_o_expo_lpi_2[3:0]),
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_270_nl = ~ data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_47_nl
      = MUX_v_4_2_2(4'b0000, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_mux_171_nl),
      (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_not_270_nl));
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_mux_171_nl = MUX_v_4_2_2(4'b1110, (FpExpoWidthDec_6U_5U_10U_1U_1U_else_FpExpoWidthDec_6U_5U_10U_1U_1U_else_and_47_nl),
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_31_nl
      = MUX_v_4_2_2((FpExpoWidthDec_6U_5U_10U_1U_1U_mux_171_nl), 4'b1111, IsNaN_6U_10U_16_land_lpi_1_dfm);
  assign or_1389_nl = or_dcpl_293 | data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1;
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_31_nl = MUX_s_1_2_2(data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_itm_6_1,
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_acc_6_svs,
      or_1389_nl);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_31_nl = MUX_s_1_2_2(data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_itm_5_1,
      data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_acc_5_svs,
      or_dcpl_293);
  assign FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_1_or_30_nl
      = ((~ (FpAdd_6U_10U_7_o_expo_lpi_2[4])) & (FpExpoWidthDec_6U_5U_10U_1U_1U_else_else_if_mux_31_nl)
      & (~ (FpExpoWidthDec_6U_5U_10U_1U_1U_else_if_mux_31_nl))) | (~ data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2)
      | IsNaN_6U_10U_16_land_lpi_1_dfm;
  assign mux_52_nl = MUX_s_1_2_2(not_tmp_81, mux_tmp_51, or_tmp_5);
  assign mux_53_nl = MUX_s_1_2_2(not_tmp_81, mux_tmp_51, or_99_cse);
  assign mux_54_nl = MUX_s_1_2_2((mux_53_nl), (mux_52_nl), nor_57_cse);
  assign mux_57_nl = MUX_s_1_2_2(not_tmp_83, mux_tmp_56, or_tmp_8);
  assign mux_58_nl = MUX_s_1_2_2(not_tmp_83, mux_tmp_56, or_109_cse);
  assign mux_59_nl = MUX_s_1_2_2((mux_58_nl), (mux_57_nl), nor_57_cse);
  assign mux_62_nl = MUX_s_1_2_2(not_tmp_85, mux_tmp_61, or_tmp_16);
  assign mux_63_nl = MUX_s_1_2_2(not_tmp_85, mux_tmp_61, or_119_cse);
  assign mux_64_nl = MUX_s_1_2_2((mux_63_nl), (mux_62_nl), nor_57_cse);
  assign mux_70_nl = MUX_s_1_2_2(not_tmp_90, mux_tmp_69, or_tmp_52);
  assign mux_71_nl = MUX_s_1_2_2(not_tmp_90, mux_tmp_69, or_134_cse);
  assign mux_72_nl = MUX_s_1_2_2((mux_71_nl), (mux_70_nl), nor_57_cse);
  assign mux_82_nl = MUX_s_1_2_2(not_tmp_96, mux_tmp_81, or_tmp_48);
  assign mux_83_nl = MUX_s_1_2_2(not_tmp_96, mux_tmp_81, or_152_cse);
  assign mux_84_nl = MUX_s_1_2_2((mux_83_nl), (mux_82_nl), nor_57_cse);
  assign mux_94_nl = MUX_s_1_2_2(not_tmp_102, mux_tmp_93, or_tmp_44);
  assign or_170_nl = nor_82_cse | IsNaN_6U_10U_6_land_1_lpi_1_dfm;
  assign mux_95_nl = MUX_s_1_2_2(not_tmp_102, mux_tmp_93, or_170_nl);
  assign mux_96_nl = MUX_s_1_2_2((mux_95_nl), (mux_94_nl), nor_57_cse);
  assign mux_107_nl = MUX_s_1_2_2(or_183_cse, or_tmp_39, nor_57_cse);
  assign and_85_nl = chn_data_in_rsci_bawt & (mux_107_nl);
  assign mux_108_nl = MUX_s_1_2_2(and_2591_cse, (and_85_nl), or_181_cse);
  assign mux_116_nl = MUX_s_1_2_2(or_196_cse, or_tmp_36, nor_57_cse);
  assign and_88_nl = chn_data_in_rsci_bawt & (mux_116_nl);
  assign mux_117_nl = MUX_s_1_2_2(and_2588_cse, (and_88_nl), or_181_cse);
  assign mux_125_nl = MUX_s_1_2_2(or_209_cse, or_tmp_33, nor_57_cse);
  assign and_91_nl = chn_data_in_rsci_bawt & (mux_125_nl);
  assign mux_126_nl = MUX_s_1_2_2(and_2585_cse, (and_91_nl), or_181_cse);
  assign mux_137_nl = MUX_s_1_2_2(or_224_cse, or_tmp_27, nor_57_cse);
  assign and_96_nl = chn_data_in_rsci_bawt & (mux_137_nl);
  assign mux_138_nl = MUX_s_1_2_2(and_2582_cse, (and_96_nl), or_181_cse);
  assign mux_146_nl = MUX_s_1_2_2(or_237_cse, or_tmp_25, nor_57_cse);
  assign and_99_nl = chn_data_in_rsci_bawt & (mux_146_nl);
  assign mux_147_nl = MUX_s_1_2_2(and_2579_cse, (and_99_nl), or_181_cse);
  assign mux_157_nl = MUX_s_1_2_2(or_256_cse, or_tmp_22, nor_57_cse);
  assign and_100_nl = chn_data_in_rsci_bawt & (mux_157_nl);
  assign mux_158_nl = MUX_s_1_2_2(and_2576_cse, (and_100_nl), or_181_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_13_nl = (~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_3)
      & and_689_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_12_nl = (~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_3)
      & and_691_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_13_nl = (~ IsNaN_6U_10U_3_land_1_lpi_1_dfm_3)
      & and_693_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_12_nl = (~ IsNaN_6U_10U_3_land_3_lpi_1_dfm_3)
      & and_695_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_13_nl = (~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_3)
      & and_697_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_12_nl = (~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_3)
      & and_699_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_13_nl = (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_3)
      & and_701_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_12_nl = (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_3)
      & and_703_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_11_nl = (~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_3)
      & and_705_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_11_nl = (~ IsNaN_6U_10U_3_land_2_lpi_1_dfm_3)
      & and_707_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_11_nl = (~ IsNaN_6U_10U_5_land_2_lpi_1_dfm_3)
      & and_709_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_11_nl = (~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_3)
      & and_711_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_nl = and_713_rgt | (IsNaN_6U_10U_1_land_lpi_1_dfm_3
      & and_715_rgt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_10_nl = (~ IsNaN_6U_10U_1_land_lpi_1_dfm_3)
      & and_715_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_nl = and_717_rgt | (IsNaN_6U_10U_3_land_lpi_1_dfm_3
      & and_719_rgt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_10_nl = (~ IsNaN_6U_10U_3_land_lpi_1_dfm_3)
      & and_719_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_or_nl = and_721_rgt | (IsNaN_6U_10U_5_land_lpi_1_dfm_3
      & and_723_rgt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_10_nl = (~ IsNaN_6U_10U_5_land_lpi_1_dfm_3)
      & and_723_rgt;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_or_nl = and_725_rgt | (IsNaN_6U_10U_7_land_lpi_1_dfm_3
      & and_727_rgt);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_10_nl = (~ IsNaN_6U_10U_7_land_lpi_1_dfm_3)
      & and_727_rgt;
  assign FpAdd_6U_10U_7_else_2_mux_8_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_7_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_6U_10U_7_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp);
  assign FpAdd_6U_10U_7_else_2_mux_9_nl = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_6U_10U_7_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp);
  assign nl_acc_16_nl = ({(~ FpAdd_6U_10U_7_if_2_and_tmp) , (FpAdd_6U_10U_7_else_2_mux_8_nl)
      , (~ FpAdd_6U_10U_7_if_2_and_tmp)}) + conv_u2u_24_25({(FpAdd_6U_10U_7_else_2_mux_9_nl)
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[24:0];
  assign FpAdd_6U_10U_7_else_2_mux_10_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_7_addend_smaller_qr_3_lpi_1_dfm_mx0),
      FpAdd_6U_10U_7_addend_larger_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_1);
  assign FpAdd_6U_10U_7_else_2_mux_11_nl = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_qr_3_lpi_1_dfm_mx0,
      FpAdd_6U_10U_7_addend_smaller_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_1);
  assign nl_acc_17_nl = ({(~ FpAdd_6U_10U_7_if_2_and_tmp_1) , (FpAdd_6U_10U_7_else_2_mux_10_nl)
      , (~ FpAdd_6U_10U_7_if_2_and_tmp_1)}) + conv_u2u_24_25({(FpAdd_6U_10U_7_else_2_mux_11_nl)
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[24:0];
  assign FpAdd_6U_10U_7_else_2_mux_12_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_7_addend_smaller_qr_2_lpi_1_dfm_mx0),
      FpAdd_6U_10U_7_addend_larger_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_2);
  assign FpAdd_6U_10U_7_else_2_mux_13_nl = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_qr_2_lpi_1_dfm_mx0,
      FpAdd_6U_10U_7_addend_smaller_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_2);
  assign nl_acc_18_nl = ({(~ FpAdd_6U_10U_7_if_2_and_tmp_2) , (FpAdd_6U_10U_7_else_2_mux_12_nl)
      , (~ FpAdd_6U_10U_7_if_2_and_tmp_2)}) + conv_u2u_24_25({(FpAdd_6U_10U_7_else_2_mux_13_nl)
      , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[24:0];
  assign FpAdd_6U_10U_7_else_2_mux_14_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_7_addend_smaller_qr_1_lpi_1_dfm_mx0),
      FpAdd_6U_10U_7_addend_larger_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_3);
  assign FpAdd_6U_10U_7_else_2_mux_15_nl = MUX_v_23_2_2(FpAdd_6U_10U_7_addend_larger_qr_1_lpi_1_dfm_mx0,
      FpAdd_6U_10U_7_addend_smaller_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_7_if_2_and_tmp_3);
  assign nl_acc_19_nl = ({(~ FpAdd_6U_10U_7_if_2_and_tmp_3) , (FpAdd_6U_10U_7_else_2_mux_14_nl)
      , (~ FpAdd_6U_10U_7_if_2_and_tmp_3)}) + conv_u2u_24_25({(FpAdd_6U_10U_7_else_2_mux_15_nl)
      , 1'b1});
  assign acc_19_nl = nl_acc_19_nl[24:0];
  assign FpAdd_6U_10U_6_else_2_mux_8_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_6_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_6U_10U_6_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp);
  assign FpAdd_6U_10U_6_else_2_mux_9_nl = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_6U_10U_6_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp);
  assign nl_acc_20_nl = ({(~ FpAdd_6U_10U_6_if_2_and_tmp) , (FpAdd_6U_10U_6_else_2_mux_8_nl)
      , (~ FpAdd_6U_10U_6_if_2_and_tmp)}) + conv_u2u_24_25({(FpAdd_6U_10U_6_else_2_mux_9_nl)
      , 1'b1});
  assign acc_20_nl = nl_acc_20_nl[24:0];
  assign FpAdd_6U_10U_6_else_2_mux_10_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_6_addend_smaller_qr_3_lpi_1_dfm_mx0),
      FpAdd_6U_10U_6_addend_larger_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_1);
  assign FpAdd_6U_10U_6_else_2_mux_11_nl = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_qr_3_lpi_1_dfm_mx0,
      FpAdd_6U_10U_6_addend_smaller_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_1);
  assign nl_acc_21_nl = ({(~ FpAdd_6U_10U_6_if_2_and_tmp_1) , (FpAdd_6U_10U_6_else_2_mux_10_nl)
      , (~ FpAdd_6U_10U_6_if_2_and_tmp_1)}) + conv_u2u_24_25({(FpAdd_6U_10U_6_else_2_mux_11_nl)
      , 1'b1});
  assign acc_21_nl = nl_acc_21_nl[24:0];
  assign FpAdd_6U_10U_6_else_2_mux_12_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_6_addend_smaller_qr_2_lpi_1_dfm_mx0),
      FpAdd_6U_10U_6_addend_larger_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_2);
  assign FpAdd_6U_10U_6_else_2_mux_13_nl = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_qr_2_lpi_1_dfm_mx0,
      FpAdd_6U_10U_6_addend_smaller_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_2);
  assign nl_acc_22_nl = ({(~ FpAdd_6U_10U_6_if_2_and_tmp_2) , (FpAdd_6U_10U_6_else_2_mux_12_nl)
      , (~ FpAdd_6U_10U_6_if_2_and_tmp_2)}) + conv_u2u_24_25({(FpAdd_6U_10U_6_else_2_mux_13_nl)
      , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[24:0];
  assign FpAdd_6U_10U_6_else_2_mux_14_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_6_addend_smaller_qr_1_lpi_1_dfm_mx0),
      FpAdd_6U_10U_6_addend_larger_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_3);
  assign FpAdd_6U_10U_6_else_2_mux_15_nl = MUX_v_23_2_2(FpAdd_6U_10U_6_addend_larger_qr_1_lpi_1_dfm_mx0,
      FpAdd_6U_10U_6_addend_smaller_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_6_if_2_and_tmp_3);
  assign nl_acc_23_nl = ({(~ FpAdd_6U_10U_6_if_2_and_tmp_3) , (FpAdd_6U_10U_6_else_2_mux_14_nl)
      , (~ FpAdd_6U_10U_6_if_2_and_tmp_3)}) + conv_u2u_24_25({(FpAdd_6U_10U_6_else_2_mux_15_nl)
      , 1'b1});
  assign acc_23_nl = nl_acc_23_nl[24:0];
  assign FpAdd_6U_10U_5_else_2_mux_8_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_5_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_6U_10U_5_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp);
  assign FpAdd_6U_10U_5_else_2_mux_9_nl = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_6U_10U_5_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp);
  assign nl_acc_24_nl = ({(~ FpAdd_6U_10U_5_if_2_and_tmp) , (FpAdd_6U_10U_5_else_2_mux_8_nl)
      , (~ FpAdd_6U_10U_5_if_2_and_tmp)}) + conv_u2u_24_25({(FpAdd_6U_10U_5_else_2_mux_9_nl)
      , 1'b1});
  assign acc_24_nl = nl_acc_24_nl[24:0];
  assign FpAdd_6U_10U_5_else_2_mux_10_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_5_addend_smaller_qr_3_lpi_1_dfm_mx0),
      FpAdd_6U_10U_5_addend_larger_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_1);
  assign FpAdd_6U_10U_5_else_2_mux_11_nl = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_qr_3_lpi_1_dfm_mx0,
      FpAdd_6U_10U_5_addend_smaller_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_1);
  assign nl_acc_25_nl = ({(~ FpAdd_6U_10U_5_if_2_and_tmp_1) , (FpAdd_6U_10U_5_else_2_mux_10_nl)
      , (~ FpAdd_6U_10U_5_if_2_and_tmp_1)}) + conv_u2u_24_25({(FpAdd_6U_10U_5_else_2_mux_11_nl)
      , 1'b1});
  assign acc_25_nl = nl_acc_25_nl[24:0];
  assign FpAdd_6U_10U_5_else_2_mux_12_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_5_addend_smaller_qr_2_lpi_1_dfm_mx0),
      FpAdd_6U_10U_5_addend_larger_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_2);
  assign FpAdd_6U_10U_5_else_2_mux_13_nl = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_qr_2_lpi_1_dfm_mx0,
      FpAdd_6U_10U_5_addend_smaller_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_2);
  assign nl_acc_26_nl = ({(~ FpAdd_6U_10U_5_if_2_and_tmp_2) , (FpAdd_6U_10U_5_else_2_mux_12_nl)
      , (~ FpAdd_6U_10U_5_if_2_and_tmp_2)}) + conv_u2u_24_25({(FpAdd_6U_10U_5_else_2_mux_13_nl)
      , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[24:0];
  assign FpAdd_6U_10U_5_else_2_mux_14_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_5_addend_smaller_qr_1_lpi_1_dfm_mx0),
      FpAdd_6U_10U_5_addend_larger_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_3);
  assign FpAdd_6U_10U_5_else_2_mux_15_nl = MUX_v_23_2_2(FpAdd_6U_10U_5_addend_larger_qr_1_lpi_1_dfm_mx0,
      FpAdd_6U_10U_5_addend_smaller_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_5_if_2_and_tmp_3);
  assign nl_acc_27_nl = ({(~ FpAdd_6U_10U_5_if_2_and_tmp_3) , (FpAdd_6U_10U_5_else_2_mux_14_nl)
      , (~ FpAdd_6U_10U_5_if_2_and_tmp_3)}) + conv_u2u_24_25({(FpAdd_6U_10U_5_else_2_mux_15_nl)
      , 1'b1});
  assign acc_27_nl = nl_acc_27_nl[24:0];
  assign FpAdd_6U_10U_4_else_2_mux_8_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_4_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_6U_10U_4_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp);
  assign FpAdd_6U_10U_4_else_2_mux_9_nl = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_6U_10U_4_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp);
  assign nl_acc_28_nl = ({(~ FpAdd_6U_10U_4_if_2_and_tmp) , (FpAdd_6U_10U_4_else_2_mux_8_nl)
      , (~ FpAdd_6U_10U_4_if_2_and_tmp)}) + conv_u2u_24_25({(FpAdd_6U_10U_4_else_2_mux_9_nl)
      , 1'b1});
  assign acc_28_nl = nl_acc_28_nl[24:0];
  assign FpAdd_6U_10U_4_else_2_mux_10_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_4_addend_smaller_qr_3_lpi_1_dfm_mx0),
      FpAdd_6U_10U_4_addend_larger_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_1);
  assign FpAdd_6U_10U_4_else_2_mux_11_nl = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_qr_3_lpi_1_dfm_mx0,
      FpAdd_6U_10U_4_addend_smaller_qr_3_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_1);
  assign nl_acc_29_nl = ({(~ FpAdd_6U_10U_4_if_2_and_tmp_1) , (FpAdd_6U_10U_4_else_2_mux_10_nl)
      , (~ FpAdd_6U_10U_4_if_2_and_tmp_1)}) + conv_u2u_24_25({(FpAdd_6U_10U_4_else_2_mux_11_nl)
      , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[24:0];
  assign FpAdd_6U_10U_4_else_2_mux_12_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_4_addend_smaller_qr_2_lpi_1_dfm_mx0),
      FpAdd_6U_10U_4_addend_larger_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_2);
  assign FpAdd_6U_10U_4_else_2_mux_13_nl = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_qr_2_lpi_1_dfm_mx0,
      FpAdd_6U_10U_4_addend_smaller_qr_2_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_2);
  assign nl_acc_30_nl = ({(~ FpAdd_6U_10U_4_if_2_and_tmp_2) , (FpAdd_6U_10U_4_else_2_mux_12_nl)
      , (~ FpAdd_6U_10U_4_if_2_and_tmp_2)}) + conv_u2u_24_25({(FpAdd_6U_10U_4_else_2_mux_13_nl)
      , 1'b1});
  assign acc_30_nl = nl_acc_30_nl[24:0];
  assign FpAdd_6U_10U_4_else_2_mux_14_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_4_addend_smaller_qr_1_lpi_1_dfm_mx0),
      FpAdd_6U_10U_4_addend_larger_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_3);
  assign FpAdd_6U_10U_4_else_2_mux_15_nl = MUX_v_23_2_2(FpAdd_6U_10U_4_addend_larger_qr_1_lpi_1_dfm_mx0,
      FpAdd_6U_10U_4_addend_smaller_qr_1_lpi_1_dfm_mx0, FpAdd_6U_10U_4_if_2_and_tmp_3);
  assign nl_acc_31_nl = ({(~ FpAdd_6U_10U_4_if_2_and_tmp_3) , (FpAdd_6U_10U_4_else_2_mux_14_nl)
      , (~ FpAdd_6U_10U_4_if_2_and_tmp_3)}) + conv_u2u_24_25({(FpAdd_6U_10U_4_else_2_mux_15_nl)
      , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[24:0];
  assign mux_209_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_311_cse);
  assign and_2562_nl = data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  assign mux_210_nl = MUX_s_1_2_2((mux_209_nl), mux_tmp_206, and_2562_nl);
  assign mux_211_nl = MUX_s_1_2_2((mux_210_nl), mux_tmp_206, IsNaN_6U_10U_16_land_12_lpi_1_dfm_3);
  assign mux_213_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_315_cse);
  assign and_2561_nl = data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_214_nl = MUX_s_1_2_2((mux_213_nl), mux_tmp_212, and_2561_nl);
  assign mux_215_nl = MUX_s_1_2_2((mux_214_nl), mux_tmp_212, IsNaN_6U_10U_16_land_8_lpi_1_dfm_3);
  assign mux_216_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_202, or_317_cse);
  assign mux_217_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_205, or_317_cse);
  assign or_316_nl = data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_3_tmp;
  assign mux_218_nl = MUX_s_1_2_2((mux_217_nl), (mux_216_nl), or_316_nl);
  assign or_319_nl = data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_220_nl = MUX_s_1_2_2(mux_tmp_219, or_tmp_303, or_319_nl);
  assign or_327_nl = data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_221_nl = MUX_s_1_2_2(mux_tmp_219, or_tmp_303, or_327_nl);
  assign mux_222_nl = MUX_s_1_2_2((mux_221_nl), (mux_220_nl), cfg_precision[1]);
  assign or_330_nl = (or_tmp_302 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_223_nl = MUX_s_1_2_2((or_330_nl), (mux_222_nl), main_stage_v_3);
  assign nor_515_nl = ~((~(and_2555_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_331_nl = (~ (cfg_precision[1])) | data_truncate_12_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_224_nl = MUX_s_1_2_2((nor_515_nl), or_tmp_303, or_331_nl);
  assign mux_225_nl = MUX_s_1_2_2(nand_147_cse, (mux_224_nl), main_stage_v_3);
  assign nand_41_nl = ~(main_stage_v_3 & (~ or_tmp_303));
  assign mux_226_nl = MUX_s_1_2_2((nand_41_nl), (mux_225_nl), nor_150_cse);
  assign mux_227_nl = MUX_s_1_2_2((mux_226_nl), (mux_223_nl), main_stage_v_2);
  assign or_336_nl = data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_229_nl = MUX_s_1_2_2(mux_tmp_228, or_tmp_320, or_336_nl);
  assign or_344_nl = data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_230_nl = MUX_s_1_2_2(mux_tmp_228, or_tmp_320, or_344_nl);
  assign mux_231_nl = MUX_s_1_2_2((mux_230_nl), (mux_229_nl), cfg_precision[1]);
  assign or_347_nl = (or_tmp_319 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_232_nl = MUX_s_1_2_2((or_347_nl), (mux_231_nl), main_stage_v_3);
  assign nor_512_nl = ~((~(and_2550_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_348_nl = (~ (cfg_precision[1])) | data_truncate_8_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_233_nl = MUX_s_1_2_2((nor_512_nl), or_tmp_320, or_348_nl);
  assign mux_234_nl = MUX_s_1_2_2(nand_147_cse, (mux_233_nl), main_stage_v_3);
  assign nand_42_nl = ~(main_stage_v_3 & (~ or_tmp_320));
  assign mux_235_nl = MUX_s_1_2_2((nand_42_nl), (mux_234_nl), nor_150_cse);
  assign mux_236_nl = MUX_s_1_2_2((mux_235_nl), (mux_232_nl), main_stage_v_2);
  assign or_353_nl = data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_238_nl = MUX_s_1_2_2(mux_tmp_237, or_tmp_337, or_353_nl);
  assign or_361_nl = data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_239_nl = MUX_s_1_2_2(mux_tmp_237, or_tmp_337, or_361_nl);
  assign mux_240_nl = MUX_s_1_2_2((mux_239_nl), (mux_238_nl), cfg_precision[1]);
  assign or_364_nl = (or_tmp_336 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_241_nl = MUX_s_1_2_2((or_364_nl), (mux_240_nl), main_stage_v_3);
  assign nor_509_nl = ~((~(and_2545_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_365_nl = (~ (cfg_precision[1])) | data_truncate_4_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_242_nl = MUX_s_1_2_2((nor_509_nl), or_tmp_337, or_365_nl);
  assign mux_243_nl = MUX_s_1_2_2(nand_147_cse, (mux_242_nl), main_stage_v_3);
  assign nand_43_nl = ~(main_stage_v_3 & (~ or_tmp_337));
  assign mux_244_nl = MUX_s_1_2_2((nand_43_nl), (mux_243_nl), nor_150_cse);
  assign mux_245_nl = MUX_s_1_2_2((mux_244_nl), (mux_241_nl), main_stage_v_2);
  assign mux_247_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_371_cse);
  assign and_2543_nl = data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_248_nl = MUX_s_1_2_2((mux_247_nl), mux_tmp_246, and_2543_nl);
  assign mux_249_nl = MUX_s_1_2_2((mux_248_nl), mux_tmp_246, IsNaN_6U_10U_16_land_11_lpi_1_dfm_3);
  assign mux_251_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_373_cse);
  assign and_2542_nl = data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2
      & data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2;
  assign mux_252_nl = MUX_s_1_2_2((mux_251_nl), mux_tmp_250, and_2542_nl);
  assign mux_253_nl = MUX_s_1_2_2((mux_252_nl), mux_tmp_250, IsNaN_6U_10U_16_land_7_lpi_1_dfm_3);
  assign mux_255_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_375_cse);
  assign and_2541_nl = data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_256_nl = MUX_s_1_2_2((mux_255_nl), mux_tmp_254, and_2541_nl);
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), mux_tmp_254, IsNaN_6U_10U_16_land_3_lpi_1_dfm_3);
  assign or_376_nl = data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_259_nl = MUX_s_1_2_2(mux_tmp_258, or_tmp_360, or_376_nl);
  assign or_384_nl = data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_260_nl = MUX_s_1_2_2(mux_tmp_258, or_tmp_360, or_384_nl);
  assign mux_261_nl = MUX_s_1_2_2((mux_260_nl), (mux_259_nl), cfg_precision[1]);
  assign or_387_nl = (or_tmp_359 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_262_nl = MUX_s_1_2_2((or_387_nl), (mux_261_nl), main_stage_v_3);
  assign nor_506_nl = ~((~(and_2537_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_388_nl = (~ (cfg_precision[1])) | data_truncate_11_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_263_nl = MUX_s_1_2_2((nor_506_nl), or_tmp_360, or_388_nl);
  assign mux_264_nl = MUX_s_1_2_2(nand_147_cse, (mux_263_nl), main_stage_v_3);
  assign nand_44_nl = ~(main_stage_v_3 & (~ or_tmp_360));
  assign mux_265_nl = MUX_s_1_2_2((nand_44_nl), (mux_264_nl), nor_150_cse);
  assign mux_266_nl = MUX_s_1_2_2((mux_265_nl), (mux_262_nl), main_stage_v_2);
  assign or_393_nl = data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_268_nl = MUX_s_1_2_2(mux_tmp_267, or_tmp_377, or_393_nl);
  assign or_401_nl = data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_269_nl = MUX_s_1_2_2(mux_tmp_267, or_tmp_377, or_401_nl);
  assign mux_270_nl = MUX_s_1_2_2((mux_269_nl), (mux_268_nl), cfg_precision[1]);
  assign or_404_nl = (or_tmp_376 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_271_nl = MUX_s_1_2_2((or_404_nl), (mux_270_nl), main_stage_v_3);
  assign nor_503_nl = ~((~(and_2532_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_405_nl = (~ (cfg_precision[1])) | data_truncate_7_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_272_nl = MUX_s_1_2_2((nor_503_nl), or_tmp_377, or_405_nl);
  assign mux_273_nl = MUX_s_1_2_2(nand_147_cse, (mux_272_nl), main_stage_v_3);
  assign nand_45_nl = ~(main_stage_v_3 & (~ or_tmp_377));
  assign mux_274_nl = MUX_s_1_2_2((nand_45_nl), (mux_273_nl), nor_150_cse);
  assign mux_275_nl = MUX_s_1_2_2((mux_274_nl), (mux_271_nl), main_stage_v_2);
  assign or_410_nl = data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_277_nl = MUX_s_1_2_2(mux_tmp_276, or_tmp_394, or_410_nl);
  assign or_418_nl = data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_278_nl = MUX_s_1_2_2(mux_tmp_276, or_tmp_394, or_418_nl);
  assign mux_279_nl = MUX_s_1_2_2((mux_278_nl), (mux_277_nl), cfg_precision[1]);
  assign or_421_nl = (or_tmp_393 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_280_nl = MUX_s_1_2_2((or_421_nl), (mux_279_nl), main_stage_v_3);
  assign nor_500_nl = ~((~(and_2527_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_422_nl = (~ (cfg_precision[1])) | data_truncate_3_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_281_nl = MUX_s_1_2_2((nor_500_nl), or_tmp_394, or_422_nl);
  assign mux_282_nl = MUX_s_1_2_2(nand_147_cse, (mux_281_nl), main_stage_v_3);
  assign nand_46_nl = ~(main_stage_v_3 & (~ or_tmp_394));
  assign mux_283_nl = MUX_s_1_2_2((nand_46_nl), (mux_282_nl), nor_150_cse);
  assign mux_284_nl = MUX_s_1_2_2((mux_283_nl), (mux_280_nl), main_stage_v_2);
  assign mux_285_nl = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_427_cse);
  assign mux_286_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_202, IsNaN_6U_10U_16_land_10_lpi_1_dfm_3);
  assign mux_287_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_205, IsNaN_6U_10U_16_land_10_lpi_1_dfm_3);
  assign mux_288_nl = MUX_s_1_2_2((mux_287_nl), (mux_286_nl), or_427_cse);
  assign and_2525_nl = data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_289_nl = MUX_s_1_2_2((mux_288_nl), (mux_285_nl), and_2525_nl);
  assign mux_290_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_202, or_429_cse);
  assign mux_292_nl = MUX_s_1_2_2(or_tmp_290, mux_tmp_291, or_181_cse);
  assign mux_293_nl = MUX_s_1_2_2(mux_tmp_201, mux_tmp_291, or_181_cse);
  assign mux_294_nl = MUX_s_1_2_2((mux_293_nl), (mux_292_nl), or_429_cse);
  assign mux_295_nl = MUX_s_1_2_2((mux_294_nl), (mux_290_nl), IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_5_tmp);
  assign mux_296_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_202, or_434_cse);
  assign mux_297_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_205, or_434_cse);
  assign or_433_nl = IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_1_tmp | data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1;
  assign mux_298_nl = MUX_s_1_2_2((mux_297_nl), (mux_296_nl), or_433_nl);
  assign or_436_nl = data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_300_nl = MUX_s_1_2_2(mux_tmp_299, or_tmp_420, or_436_nl);
  assign or_444_nl = data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_301_nl = MUX_s_1_2_2(mux_tmp_299, or_tmp_420, or_444_nl);
  assign mux_302_nl = MUX_s_1_2_2((mux_301_nl), (mux_300_nl), cfg_precision[1]);
  assign or_447_nl = (or_tmp_419 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_303_nl = MUX_s_1_2_2((or_447_nl), (mux_302_nl), main_stage_v_3);
  assign nor_497_nl = ~((~(and_2517_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_448_nl = (~ (cfg_precision[1])) | data_truncate_10_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_304_nl = MUX_s_1_2_2((nor_497_nl), or_tmp_420, or_448_nl);
  assign mux_305_nl = MUX_s_1_2_2(nand_147_cse, (mux_304_nl), main_stage_v_3);
  assign nand_47_nl = ~(main_stage_v_3 & (~ or_tmp_420));
  assign mux_306_nl = MUX_s_1_2_2((nand_47_nl), (mux_305_nl), nor_150_cse);
  assign mux_307_nl = MUX_s_1_2_2((mux_306_nl), (mux_303_nl), main_stage_v_2);
  assign mux_314_nl = MUX_s_1_2_2(or_tmp_438, mux_tmp_313, or_181_cse);
  assign mux_315_nl = MUX_s_1_2_2(or_tmp_290, mux_tmp_313, or_181_cse);
  assign mux_316_nl = MUX_s_1_2_2((mux_315_nl), (mux_314_nl), data_truncate_6_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_458_nl = data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_318_nl = MUX_s_1_2_2(mux_tmp_317, or_tmp_442, or_458_nl);
  assign or_466_nl = data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_319_nl = MUX_s_1_2_2(mux_tmp_317, or_tmp_442, or_466_nl);
  assign mux_320_nl = MUX_s_1_2_2((mux_319_nl), (mux_318_nl), cfg_precision[1]);
  assign or_469_nl = (or_tmp_441 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_321_nl = MUX_s_1_2_2((or_469_nl), (mux_320_nl), main_stage_v_3);
  assign nor_494_nl = ~((~(and_2512_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_470_nl = (~ (cfg_precision[1])) | data_truncate_2_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_322_nl = MUX_s_1_2_2((nor_494_nl), or_tmp_442, or_470_nl);
  assign mux_323_nl = MUX_s_1_2_2(nand_147_cse, (mux_322_nl), main_stage_v_3);
  assign nand_48_nl = ~(main_stage_v_3 & (~ or_tmp_442));
  assign mux_324_nl = MUX_s_1_2_2((nand_48_nl), (mux_323_nl), nor_150_cse);
  assign mux_325_nl = MUX_s_1_2_2((mux_324_nl), (mux_321_nl), main_stage_v_2);
  assign mux_326_nl = MUX_s_1_2_2(mux_tmp_205, mux_tmp_202, or_476_cse);
  assign mux_327_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_476_cse);
  assign or_475_nl = (data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | IsNaN_6U_10U_16_land_9_lpi_1_dfm_3;
  assign mux_328_nl = MUX_s_1_2_2((mux_327_nl), (mux_326_nl), or_475_nl);
  assign mux_330_nl = MUX_s_1_2_2(or_tmp_290, mux_tmp_329, or_181_cse);
  assign mux_331_nl = MUX_s_1_2_2((mux_330_nl), mux_tmp_202, IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_4_tmp);
  assign mux_332_nl = MUX_s_1_2_2(mux_tmp_201, mux_tmp_329, or_181_cse);
  assign mux_333_nl = MUX_s_1_2_2((mux_332_nl), mux_tmp_207, IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_4_tmp);
  assign or_478_nl = (data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | IsNaN_6U_10U_16_land_5_lpi_1_dfm_3;
  assign mux_334_nl = MUX_s_1_2_2((mux_333_nl), (mux_331_nl), or_478_nl);
  assign mux_335_nl = MUX_s_1_2_2(mux_tmp_207, mux_tmp_202, and_2507_cse);
  assign mux_336_nl = MUX_s_1_2_2((mux_335_nl), mux_tmp_202, IsNaN_6U_10U_16_land_1_lpi_1_dfm_3);
  assign mux_337_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_205, and_2507_cse);
  assign mux_338_nl = MUX_s_1_2_2((mux_337_nl), mux_tmp_205, IsNaN_6U_10U_16_land_1_lpi_1_dfm_3);
  assign or_481_nl = data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      IsNaN_6U_10U_16_IsNaN_6U_10U_16_nor_tmp;
  assign mux_339_nl = MUX_s_1_2_2((mux_338_nl), (mux_336_nl), or_481_nl);
  assign or_482_nl = data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_341_nl = MUX_s_1_2_2(mux_tmp_340, or_tmp_466, or_482_nl);
  assign or_490_nl = data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_342_nl = MUX_s_1_2_2(mux_tmp_340, or_tmp_466, or_490_nl);
  assign mux_343_nl = MUX_s_1_2_2((mux_342_nl), (mux_341_nl), cfg_precision[1]);
  assign or_493_nl = (or_tmp_465 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_344_nl = MUX_s_1_2_2((or_493_nl), (mux_343_nl), main_stage_v_3);
  assign nor_491_nl = ~((~(and_2503_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_494_nl = (~ (cfg_precision[1])) | data_truncate_9_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_345_nl = MUX_s_1_2_2((nor_491_nl), or_tmp_466, or_494_nl);
  assign mux_346_nl = MUX_s_1_2_2(nand_147_cse, (mux_345_nl), main_stage_v_3);
  assign nand_49_nl = ~(main_stage_v_3 & (~ or_tmp_466));
  assign mux_347_nl = MUX_s_1_2_2((nand_49_nl), (mux_346_nl), nor_150_cse);
  assign mux_348_nl = MUX_s_1_2_2((mux_347_nl), (mux_344_nl), main_stage_v_2);
  assign mux_352_nl = MUX_s_1_2_2(or_tmp_438, mux_tmp_351, or_181_cse);
  assign mux_353_nl = MUX_s_1_2_2(or_tmp_290, mux_tmp_351, or_181_cse);
  assign mux_354_nl = MUX_s_1_2_2((mux_353_nl), (mux_352_nl), data_truncate_5_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2);
  assign or_502_nl = data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1 |
      data_truncate_nor_tmp_4;
  assign mux_356_nl = MUX_s_1_2_2(mux_tmp_355, or_tmp_486, or_502_nl);
  assign or_510_nl = data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_357_nl = MUX_s_1_2_2(mux_tmp_355, or_tmp_486, or_510_nl);
  assign mux_358_nl = MUX_s_1_2_2((mux_357_nl), (mux_356_nl), cfg_precision[1]);
  assign or_513_nl = (or_tmp_485 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_359_nl = MUX_s_1_2_2((or_513_nl), (mux_358_nl), main_stage_v_3);
  assign nor_488_nl = ~((~(and_2498_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_514_nl = (~ (cfg_precision[1])) | data_truncate_1_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_360_nl = MUX_s_1_2_2((nor_488_nl), or_tmp_486, or_514_nl);
  assign mux_361_nl = MUX_s_1_2_2(nand_147_cse, (mux_360_nl), main_stage_v_3);
  assign nand_50_nl = ~(main_stage_v_3 & (~ or_tmp_486));
  assign mux_362_nl = MUX_s_1_2_2((nand_50_nl), (mux_361_nl), nor_150_cse);
  assign mux_363_nl = MUX_s_1_2_2((mux_362_nl), (mux_359_nl), main_stage_v_2);
  assign or_522_nl = (~(IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_tmp | IsNaN_6U_10U_16_nor_15_tmp
      | (~ data_truncate_nor_tmp_4) | (~ main_stage_v_3))) | mux_tmp_364;
  assign mux_365_nl = MUX_s_1_2_2((or_522_nl), or_521_cse, data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_525_nl = (data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      & data_truncate_nor_tmp_4 & main_stage_v_3) | m_row0_unequal_tmp_3 | (~ main_stage_v_2);
  assign or_523_nl = IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_15_itm | IsNaN_6U_10U_16_nor_15_itm;
  assign mux_366_nl = MUX_s_1_2_2(or_527_cse, (or_525_nl), or_523_nl);
  assign mux_367_nl = MUX_s_1_2_2((mux_366_nl), (mux_365_nl), cfg_precision[1]);
  assign or_529_nl = (data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | (~(or_tmp_510 & (~ mux_tmp_201)));
  assign mux_369_nl = MUX_s_1_2_2(mux_tmp_201, (or_529_nl), and_2495_cse);
  assign mux_370_nl = MUX_s_1_2_2((mux_369_nl), (mux_367_nl), or_181_cse);
  assign or_530_nl = data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_372_nl = MUX_s_1_2_2(mux_tmp_371, or_tmp_514, or_530_nl);
  assign or_538_nl = data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_373_nl = MUX_s_1_2_2(mux_tmp_371, or_tmp_514, or_538_nl);
  assign mux_374_nl = MUX_s_1_2_2((mux_373_nl), (mux_372_nl), cfg_precision[1]);
  assign or_541_nl = (or_tmp_513 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_375_nl = MUX_s_1_2_2((or_541_nl), (mux_374_nl), main_stage_v_3);
  assign nor_485_nl = ~((~(and_2487_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_542_nl = (~ (cfg_precision[1])) | data_truncate_16_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_376_nl = MUX_s_1_2_2((nor_485_nl), or_tmp_514, or_542_nl);
  assign mux_377_nl = MUX_s_1_2_2(nand_147_cse, (mux_376_nl), main_stage_v_3);
  assign nand_52_nl = ~(main_stage_v_3 & (~ or_tmp_514));
  assign mux_378_nl = MUX_s_1_2_2((nand_52_nl), (mux_377_nl), nor_150_cse);
  assign mux_379_nl = MUX_s_1_2_2((mux_378_nl), (mux_375_nl), main_stage_v_2);
  assign mux_381_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_548_cse);
  assign and_2485_nl = data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_382_nl = MUX_s_1_2_2((mux_381_nl), mux_tmp_380, and_2485_nl);
  assign mux_383_nl = MUX_s_1_2_2((mux_382_nl), mux_tmp_380, IsNaN_6U_10U_16_land_15_lpi_1_dfm_3);
  assign or_549_nl = data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_385_nl = MUX_s_1_2_2(mux_tmp_384, or_tmp_533, or_549_nl);
  assign or_557_nl = data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_386_nl = MUX_s_1_2_2(mux_tmp_384, or_tmp_533, or_557_nl);
  assign mux_387_nl = MUX_s_1_2_2((mux_386_nl), (mux_385_nl), cfg_precision[1]);
  assign or_560_nl = (or_tmp_532 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_388_nl = MUX_s_1_2_2((or_560_nl), (mux_387_nl), main_stage_v_3);
  assign nor_482_nl = ~((~(and_2481_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_561_nl = (~ (cfg_precision[1])) | data_truncate_15_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_389_nl = MUX_s_1_2_2((nor_482_nl), or_tmp_533, or_561_nl);
  assign mux_390_nl = MUX_s_1_2_2(nand_147_cse, (mux_389_nl), main_stage_v_3);
  assign nand_53_nl = ~(main_stage_v_3 & (~ or_tmp_533));
  assign mux_391_nl = MUX_s_1_2_2((nand_53_nl), (mux_390_nl), nor_150_cse);
  assign mux_392_nl = MUX_s_1_2_2((mux_391_nl), (mux_388_nl), main_stage_v_2);
  assign mux_394_nl = MUX_s_1_2_2(mux_tmp_208, mux_tmp_207, or_567_cse);
  assign and_2479_nl = data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2;
  assign mux_395_nl = MUX_s_1_2_2((mux_394_nl), mux_tmp_393, and_2479_nl);
  assign mux_396_nl = MUX_s_1_2_2((mux_395_nl), mux_tmp_393, IsNaN_6U_10U_16_land_14_lpi_1_dfm_3);
  assign or_568_nl = data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_398_nl = MUX_s_1_2_2(mux_tmp_397, or_tmp_552, or_568_nl);
  assign or_576_nl = data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_399_nl = MUX_s_1_2_2(mux_tmp_397, or_tmp_552, or_576_nl);
  assign mux_400_nl = MUX_s_1_2_2((mux_399_nl), (mux_398_nl), cfg_precision[1]);
  assign or_579_nl = (or_tmp_551 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_401_nl = MUX_s_1_2_2((or_579_nl), (mux_400_nl), main_stage_v_3);
  assign nor_479_nl = ~((~(and_2475_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_580_nl = (~ (cfg_precision[1])) | data_truncate_14_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_402_nl = MUX_s_1_2_2((nor_479_nl), or_tmp_552, or_580_nl);
  assign mux_403_nl = MUX_s_1_2_2(nand_147_cse, (mux_402_nl), main_stage_v_3);
  assign nand_54_nl = ~(main_stage_v_3 & (~ or_tmp_552));
  assign mux_404_nl = MUX_s_1_2_2((nand_54_nl), (mux_403_nl), nor_150_cse);
  assign mux_405_nl = MUX_s_1_2_2((mux_404_nl), (mux_401_nl), main_stage_v_2);
  assign or_588_nl = (~(IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_tmp | IsNaN_6U_10U_16_nor_12_tmp
      | (~ data_truncate_nor_tmp_4) | (~ main_stage_v_3))) | mux_tmp_364;
  assign mux_407_nl = MUX_s_1_2_2((or_588_nl), or_521_cse, data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1);
  assign or_591_nl = (data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      & data_truncate_nor_tmp_4 & main_stage_v_3) | m_row0_unequal_tmp_3 | (~ main_stage_v_2);
  assign or_589_nl = IsNaN_6U_10U_16_IsNaN_6U_10U_16_nand_12_itm | IsNaN_6U_10U_16_nor_12_itm;
  assign mux_408_nl = MUX_s_1_2_2(or_527_cse, (or_591_nl), or_589_nl);
  assign mux_409_nl = MUX_s_1_2_2((mux_408_nl), (mux_407_nl), cfg_precision[1]);
  assign or_595_nl = (data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_2
      & data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st_2)
      | (~(or_tmp_576 & (~ mux_tmp_201)));
  assign mux_411_nl = MUX_s_1_2_2(mux_tmp_201, (or_595_nl), and_2495_cse);
  assign mux_412_nl = MUX_s_1_2_2((mux_411_nl), (mux_409_nl), or_181_cse);
  assign or_596_nl = data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_414_nl = MUX_s_1_2_2(mux_tmp_413, or_tmp_580, or_596_nl);
  assign or_604_nl = data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_if_slc_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_6_svs_st
      | data_truncate_nor_tmp_4;
  assign mux_415_nl = MUX_s_1_2_2(mux_tmp_413, or_tmp_580, or_604_nl);
  assign mux_416_nl = MUX_s_1_2_2((mux_415_nl), (mux_414_nl), cfg_precision[1]);
  assign or_607_nl = (or_tmp_579 & main_stage_v_4 & reg_chn_data_out_rsci_ld_core_psct_cse
      & (~ chn_data_out_rsci_bawt)) | m_row0_unequal_tmp_3;
  assign mux_417_nl = MUX_s_1_2_2((or_607_nl), (mux_416_nl), main_stage_v_3);
  assign nor_476_nl = ~((~(and_2464_cse | m_row0_unequal_tmp_4)) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt);
  assign or_608_nl = (~ (cfg_precision[1])) | data_truncate_13_FpExpoWidthDec_6U_5U_10U_1U_1U_acc_itm_6_1
      | data_truncate_nor_tmp_4;
  assign mux_418_nl = MUX_s_1_2_2((nor_476_nl), or_tmp_580, or_608_nl);
  assign mux_419_nl = MUX_s_1_2_2(nand_147_cse, (mux_418_nl), main_stage_v_3);
  assign nand_56_nl = ~(main_stage_v_3 & (~ or_tmp_580));
  assign mux_420_nl = MUX_s_1_2_2((nand_56_nl), (mux_419_nl), nor_150_cse);
  assign mux_421_nl = MUX_s_1_2_2((mux_420_nl), (mux_417_nl), main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_6_o_mant_and_8_nl = (~ IsNaN_6U_10U_7_land_lpi_1_dfm_3)
      & FpAdd_6U_10U_3_o_mant_lpi_1_dfm_2_mx0c1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_4_o_mant_and_8_nl = (~ IsNaN_6U_10U_5_land_lpi_1_dfm_3)
      & FpAdd_6U_10U_2_o_mant_lpi_1_dfm_2_mx0c1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_8_nl = (~ IsNaN_6U_10U_3_land_lpi_1_dfm_3)
      & FpAdd_6U_10U_1_o_mant_lpi_1_dfm_2_mx0c1;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_nl = (~ IsNaN_6U_10U_1_land_lpi_1_dfm_3)
      & FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0c1;
  assign nor_3_nl = ~(nor_562_cse | (cfg_precision!=2'b10) | (~ chn_data_in_rsci_bawt));
  assign mux_2_nl = MUX_s_1_2_2(or_109_cse, or_tmp_8, nor_3_nl);
  assign nand_9_nl = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2615_nl = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_14_nl = MUX_s_1_2_2((and_2615_nl), (nand_9_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm);
  assign nand_13_nl = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2613_nl = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_1_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_17_nl = MUX_s_1_2_2((and_2613_nl), (nand_13_nl), IsNaN_6U_10U_2_land_2_lpi_1_dfm);
  assign mux_19_nl = MUX_s_1_2_2((~ nand_tmp_16), nand_tmp_15, IsNaN_6U_10U_3_land_3_lpi_1_dfm);
  assign mux_21_nl = MUX_s_1_2_2((mux_19_nl), nand_tmp_15, IsNaN_6U_10U_2_land_3_lpi_1_dfm);
  assign nand_17_nl = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2612_nl = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_2_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_22_nl = MUX_s_1_2_2((and_2612_nl), (nand_17_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm);
  assign mux_23_nl = MUX_s_1_2_2((~ nand_tmp_16), nand_tmp_15, or_224_cse);
  assign mux_36_nl = MUX_s_1_2_2(mux_tmp_35, nand_tmp_31, nor_82_cse);
  assign mux_37_nl = MUX_s_1_2_2(mux_tmp_35, nand_tmp_31, IsNaN_6U_10U_7_land_1_lpi_1_dfm);
  assign or_48_nl = (~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp;
  assign mux_38_nl = MUX_s_1_2_2(and_tmp_1, or_tmp_45, or_48_nl);
  assign nand_32_nl = ~((~((~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35);
  assign mux_39_nl = MUX_s_1_2_2((nand_32_nl), (mux_38_nl), IsNaN_6U_10U_7_land_1_lpi_1_dfm);
  assign and_2604_nl = (~((~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35;
  assign nand_151_nl = ~(((~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_1_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_1_tmp)
      & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_52_nl = (~ IsNaN_6U_10U_7_land_2_lpi_1_dfm) | IsNaN_6U_10U_6_land_2_lpi_1_dfm;
  assign mux_42_nl = MUX_s_1_2_2((nand_151_nl), (and_2604_nl), or_52_nl);
  assign or_56_nl = nor_70_cse | IsNaN_6U_10U_6_land_3_lpi_1_dfm | and_dcpl_52;
  assign and_74_nl = or_134_cse & nand_tmp_2;
  assign mux_43_nl = MUX_s_1_2_2((and_74_nl), (or_56_nl), or_tmp_52);
  assign or_60_nl = or_tmp_57 | and_dcpl_52;
  assign and_75_nl = or_tmp_57 & nand_tmp_2;
  assign mux_44_nl = MUX_s_1_2_2((and_75_nl), (or_60_nl), or_tmp_52);
  assign nor_561_nl = ~((~ IsNaN_6U_10U_7_land_3_lpi_1_dfm) | IsNaN_6U_10U_6_land_3_lpi_1_dfm
      | and_dcpl_52);
  assign nand_150_nl = ~(((~ IsNaN_6U_10U_7_land_3_lpi_1_dfm) | IsNaN_6U_10U_6_land_3_lpi_1_dfm)
      & nand_tmp_2);
  assign or_62_nl = (~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_2_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_2_tmp;
  assign mux_45_nl = MUX_s_1_2_2((nand_150_nl), (nor_561_nl), or_62_nl);
  assign mux_431_nl = MUX_s_1_2_2(not_tmp_203, mux_tmp_429, or_tmp_19);
  assign mux_432_nl = MUX_s_1_2_2(not_tmp_203, mux_tmp_429, or_623_cse);
  assign mux_433_nl = MUX_s_1_2_2((mux_432_nl), (mux_431_nl), nor_57_cse);
  assign mux_434_nl = MUX_s_1_2_2(not_tmp_203, (mux_433_nl), chn_data_in_rsci_bawt);
  assign mux_437_nl = MUX_s_1_2_2(not_tmp_204, mux_tmp_435, or_tmp_65);
  assign mux_438_nl = MUX_s_1_2_2(not_tmp_204, mux_tmp_435, or_629_cse);
  assign mux_439_nl = MUX_s_1_2_2((mux_438_nl), (mux_437_nl), nor_57_cse);
  assign mux_440_nl = MUX_s_1_2_2(not_tmp_204, (mux_439_nl), chn_data_in_rsci_bawt);
  assign mux_444_nl = MUX_s_1_2_2(or_638_cse, or_tmp_42, nor_57_cse);
  assign and_126_nl = chn_data_in_rsci_bawt & (mux_444_nl);
  assign and_2632_nl = IsNaN_6U_10U_5_land_lpi_1_dfm_3 & main_stage_v_1;
  assign mux_445_nl = MUX_s_1_2_2((and_2632_nl), main_stage_v_1, IsNaN_6U_10U_4_land_lpi_1_dfm_st_2);
  assign mux_446_nl = MUX_s_1_2_2((mux_445_nl), (and_126_nl), or_181_cse);
  assign mux_451_nl = MUX_s_1_2_2(or_648_cse, or_tmp_30, nor_57_cse);
  assign and_127_nl = chn_data_in_rsci_bawt & (mux_451_nl);
  assign and_2633_nl = IsNaN_6U_10U_3_land_lpi_1_dfm_3 & main_stage_v_1;
  assign mux_452_nl = MUX_s_1_2_2((and_2633_nl), main_stage_v_1, IsNaN_6U_10U_2_land_lpi_1_dfm_st_2);
  assign mux_453_nl = MUX_s_1_2_2((mux_452_nl), (and_127_nl), or_181_cse);
  assign data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_sva));
  assign data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_1[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_15_sva));
  assign data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_2[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_14_sva));
  assign data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_3[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_13_sva));
  assign data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_4[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_12_sva));
  assign data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_5[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_11_sva));
  assign data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_6[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_10_sva));
  assign data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_7[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_9_sva));
  assign data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_8[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_8_sva));
  assign data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_9[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_7_sva));
  assign data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_10[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_6_sva));
  assign data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_11[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_5_sva));
  assign data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_12[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_4_sva));
  assign data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_13[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_3_sva));
  assign data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_14[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_2_sva));
  assign data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_nor_2_nl = ~(MUX_v_6_2_2((z_out_15[6:1]),
      6'b111111, IntShiftRight_18U_2U_8U_obits_fixed_nor_ovfl_1_sva));
  assign data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva));
  assign data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva));
  assign data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_sva));
  assign data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_15[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva));
  assign data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_15[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva));
  assign data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_15[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_15_sva));
  assign data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_14[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva));
  assign data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_14[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva));
  assign data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_14[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_14_sva));
  assign data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_13[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva));
  assign data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_13[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva));
  assign data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_13[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_13_sva));
  assign data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_12[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva));
  assign data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_12[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva));
  assign data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_12[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_12_sva));
  assign data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_11[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva));
  assign data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_11[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva));
  assign data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_11[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_11_sva));
  assign data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_10[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva));
  assign data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_10[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva));
  assign data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_10[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_10_sva));
  assign data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_9[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva));
  assign data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_9[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva));
  assign data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_9[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_9_sva));
  assign data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_8[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva));
  assign data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_8[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva));
  assign data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_8[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_8_sva));
  assign data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_7[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva));
  assign data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_7[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva));
  assign data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_7[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_7_sva));
  assign data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_6[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva));
  assign data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_6[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva));
  assign data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_6[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_6_sva));
  assign data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_5[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva));
  assign data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_5[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva));
  assign data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_5[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_5_sva));
  assign data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_4[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva));
  assign data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_4[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva));
  assign data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_4[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_4_sva));
  assign data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_3[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva));
  assign data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_3[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva));
  assign data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_3[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_3_sva));
  assign data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_2[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva));
  assign data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_2[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva));
  assign data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_2[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_2_sva));
  assign data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_5_nl = ~(MUX_v_6_2_2((z_out_1[6:1]),
      6'b111111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva));
  assign data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_4_nl = ~(MUX_v_4_2_2((z_out_1[13:10]),
      4'b1111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva));
  assign data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_nor_2_nl = ~(MUX_v_3_2_2((z_out_1[9:7]),
      3'b111, IntShiftRight_18U_2U_16U_obits_fixed_nor_ovfl_1_sva));
  assign and_2638_nl = (~((~ main_stage_v_3) | m_row0_unequal_tmp_4)) & IsNaN_6U_10U_9_land_1_lpi_1_dfm_5;
  assign mux_544_nl = MUX_s_1_2_2((and_2638_nl), nor_439_cse, or_181_cse);
  assign and_2624_nl = or_tmp_723 & or_tmp_721;
  assign mux_545_nl = MUX_s_1_2_2(or_tmp_721, (and_2624_nl), cfg_precision[1]);
  assign mux_546_nl = MUX_s_1_2_2((mux_545_nl), or_tmp_721, cfg_precision[0]);
  assign or_738_nl = IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_3 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign mux_547_nl = MUX_s_1_2_2((mux_546_nl), or_tmp_721, or_738_nl);
  assign nor_434_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | ((~ IsNaN_6U_10U_12_land_2_lpi_1_dfm_4)
      & (mux_547_nl)));
  assign nor_436_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_11_land_2_lpi_1_dfm_5
      | (~(IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_3))))));
  assign mux_549_nl = MUX_s_1_2_2((nor_436_nl), (nor_434_nl), or_181_cse);
  assign and_2622_nl = or_tmp_738 & or_tmp_736;
  assign mux_550_nl = MUX_s_1_2_2(or_tmp_736, (and_2622_nl), cfg_precision[1]);
  assign mux_551_nl = MUX_s_1_2_2((mux_550_nl), or_tmp_736, cfg_precision[0]);
  assign or_753_nl = IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_3 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign mux_552_nl = MUX_s_1_2_2((mux_551_nl), or_tmp_736, or_753_nl);
  assign nor_429_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | ((~ IsNaN_6U_10U_12_land_3_lpi_1_dfm_4)
      & (mux_552_nl)));
  assign nor_431_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_11_land_3_lpi_1_dfm_5
      | (~(IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_5
      | (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_3))))));
  assign mux_554_nl = MUX_s_1_2_2((nor_431_nl), (nor_429_nl), or_181_cse);
  assign and_2620_nl = or_tmp_753 & or_tmp_751;
  assign mux_555_nl = MUX_s_1_2_2(or_tmp_751, (and_2620_nl), cfg_precision[1]);
  assign mux_556_nl = MUX_s_1_2_2((mux_555_nl), or_tmp_751, cfg_precision[0]);
  assign or_768_nl = IsNaN_6U_10U_8_land_lpi_1_dfm_st_3 | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign mux_557_nl = MUX_s_1_2_2((mux_556_nl), or_tmp_751, or_768_nl);
  assign nor_424_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3 | ((~ IsNaN_6U_10U_12_land_lpi_1_dfm_4)
      & (mux_557_nl)));
  assign nor_426_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_11_land_lpi_1_dfm_5
      | (~(IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 | IsNaN_6U_10U_8_land_lpi_1_dfm_5 |
      (~ IsNaN_6U_10U_9_land_lpi_1_dfm_3))))));
  assign mux_559_nl = MUX_s_1_2_2((nor_426_nl), (nor_424_nl), or_181_cse);
  assign nor_418_nl = ~((~((~(IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_1_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_1_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_1_lpi_1_dfm_st)) | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign nor_421_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_14_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_1_lpi_1_dfm_5 | (~(IsNaN_6U_10U_12_land_1_lpi_1_dfm_st_4
      | IsNaN_6U_10U_9_land_1_lpi_1_dfm_5 | (~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_5))))));
  assign mux_560_nl = MUX_s_1_2_2((nor_421_nl), (nor_418_nl), or_181_cse);
  assign nor_413_nl = ~((~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign or_795_nl = IsNaN_6U_10U_13_nor_1_itm_2 | IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign mux_561_nl = MUX_s_1_2_2(or_796_cse, (or_795_nl), nor_57_cse);
  assign nor_414_nl = ~(IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3 | IsNaN_6U_10U_12_land_2_lpi_1_dfm_4
      | (mux_561_nl));
  assign mux_562_nl = MUX_s_1_2_2((nor_414_nl), (nor_413_nl), or_tmp_774);
  assign nor_415_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_14_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_2_lpi_1_dfm_5 | (~(IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_4
      | IsNaN_6U_10U_11_land_2_lpi_1_dfm_5 | (~ IsNaN_6U_10U_13_land_2_lpi_1_dfm_3))))));
  assign mux_563_nl = MUX_s_1_2_2((nor_415_nl), (mux_562_nl), or_181_cse);
  assign nor_407_nl = ~((~((~(IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_3_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_3_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st)) | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign nor_410_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_14_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_3_lpi_1_dfm_5 | (~(IsNaN_6U_10U_12_land_3_lpi_1_dfm_st_4
      | IsNaN_6U_10U_11_land_3_lpi_1_dfm_5 | (~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_5))))));
  assign mux_564_nl = MUX_s_1_2_2((nor_410_nl), (nor_407_nl), or_181_cse);
  assign nor_401_nl = ~((~((~(IsNaN_6U_10U_12_land_lpi_1_dfm_st_3 | (~ IsNaN_6U_10U_13_land_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_lpi_1_dfm_4)) | IsNaN_6U_10U_10_land_lpi_1_dfm_4 | IsNaN_6U_10U_14_land_lpi_1_dfm_st))
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3);
  assign nor_404_nl = ~((~ main_stage_v_3) | m_row0_unequal_tmp_4 | (~(IsNaN_6U_10U_14_land_lpi_1_dfm_5
      | IsNaN_6U_10U_10_land_lpi_1_dfm_5 | (~(IsNaN_6U_10U_12_land_lpi_1_dfm_st_4
      | IsNaN_6U_10U_11_land_lpi_1_dfm_5 | (~ IsNaN_6U_10U_13_land_lpi_1_dfm_5))))));
  assign mux_565_nl = MUX_s_1_2_2((nor_404_nl), (nor_401_nl), or_181_cse);
  assign nor_399_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_10_land_1_lpi_1_dfm_st_3
      | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_1_lpi_1_dfm_st);
  assign nor_400_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_14_land_1_lpi_1_dfm_st_4
      | m_row0_unequal_tmp_4 | IsNaN_6U_10U_14_land_1_lpi_1_dfm_5 | (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_5));
  assign mux_566_nl = MUX_s_1_2_2((nor_400_nl), (nor_399_nl), or_181_cse);
  assign nor_397_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_10_land_2_lpi_1_dfm_st_3
      | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st);
  assign nor_398_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st_4
      | m_row0_unequal_tmp_4 | IsNaN_6U_10U_14_land_2_lpi_1_dfm_5 | (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_5));
  assign mux_567_nl = MUX_s_1_2_2((nor_398_nl), (nor_397_nl), or_181_cse);
  assign nor_395_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_10_land_3_lpi_1_dfm_st_3
      | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st);
  assign nor_396_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st_4
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_5 | m_row0_unequal_tmp_4 | (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_5));
  assign mux_568_nl = MUX_s_1_2_2((nor_396_nl), (nor_395_nl), or_181_cse);
  assign nor_393_nl = ~((~ main_stage_v_2) | IsNaN_6U_10U_10_land_lpi_1_dfm_st_3
      | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_15_land_lpi_1_dfm_4) | IsNaN_6U_10U_14_land_lpi_1_dfm_st);
  assign nor_394_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_14_land_lpi_1_dfm_st_4
      | m_row0_unequal_tmp_4 | IsNaN_6U_10U_14_land_lpi_1_dfm_5 | (~ IsNaN_6U_10U_15_land_lpi_1_dfm_5));
  assign mux_569_nl = MUX_s_1_2_2((nor_394_nl), (nor_393_nl), or_181_cse);
  assign mux_604_nl = MUX_s_1_2_2(mux_tmp_603, or_tmp_923, IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp);
  assign mux_605_nl = MUX_s_1_2_2(mux_tmp_603, or_tmp_923, IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp);
  assign mux_606_nl = MUX_s_1_2_2(mux_tmp_603, or_tmp_923, IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp);
  assign nand_21_nl = ~((~(IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp | (~ chn_data_in_rsci_bawt)))
      & not_tmp_35);
  assign and_2610_nl = IsNaN_6U_10U_2_IsNaN_6U_10U_2_and_3_tmp & chn_data_in_rsci_bawt
      & not_tmp_35;
  assign mux_25_nl = MUX_s_1_2_2((and_2610_nl), (nand_21_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_st);
  assign and_2602_nl = (~((~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp
      | (~ chn_data_in_rsci_bawt))) & not_tmp_35;
  assign nand_149_nl = ~(((~ IsNaN_6U_10U_7_IsNaN_6U_10U_7_and_3_tmp) | IsNaN_6U_10U_6_IsNaN_6U_10U_6_and_3_tmp)
      & chn_data_in_rsci_bawt & not_tmp_35);
  assign or_69_nl = (~ IsNaN_6U_10U_7_land_lpi_1_dfm) | IsNaN_6U_10U_6_land_lpi_1_dfm_st;
  assign mux_48_nl = MUX_s_1_2_2((nand_149_nl), (and_2602_nl), or_69_nl);
  assign or_944_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | (~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp)
      | IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nand_1_tmp
      | IsNaN_6U_10U_10_nor_1_tmp;
  assign or_945_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_10_land_2_lpi_1_dfm_4) | IsNaN_6U_10U_12_land_2_lpi_1_dfm_4;
  assign or_946_nl = IsNaN_6U_10U_13_nor_1_itm_2 | IsNaN_6U_10U_13_IsNaN_6U_10U_13_nand_1_itm_2
      | (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_10_land_2_lpi_1_dfm_4) | IsNaN_6U_10U_12_land_2_lpi_1_dfm_4;
  assign mux_609_nl = MUX_s_1_2_2((or_946_nl), (or_945_nl), IsNaN_6U_10U_12_land_2_lpi_1_dfm_st_3);
  assign mux_610_nl = MUX_s_1_2_2((mux_609_nl), (or_944_nl), or_181_cse);
  assign or_948_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp
      | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_1_tmp | IsNaN_6U_10U_9_nor_1_tmp;
  assign or_951_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4
      | or_tmp_723;
  assign mux_612_nl = MUX_s_1_2_2((or_951_nl), (or_948_nl), or_181_cse);
  assign or_953_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | (~ IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp)
      | (~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp) | IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp;
  assign or_954_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_13_land_3_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_4) | (~ IsNaN_6U_10U_10_land_3_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_3_lpi_1_dfm_4;
  assign mux_613_nl = MUX_s_1_2_2((or_954_nl), (or_953_nl), or_181_cse);
  assign or_956_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp
      | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_2_tmp | IsNaN_6U_10U_9_nor_2_tmp;
  assign or_959_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4
      | or_tmp_738;
  assign mux_615_nl = MUX_s_1_2_2((or_959_nl), (or_956_nl), or_181_cse);
  assign or_961_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | (~ IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp)
      | (~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp) | IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp;
  assign or_962_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_13_land_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_8_land_lpi_1_dfm_4) | (~ IsNaN_6U_10U_10_land_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_lpi_1_dfm_4;
  assign mux_616_nl = MUX_s_1_2_2((or_962_nl), (or_961_nl), or_181_cse);
  assign or_964_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp
      | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nand_3_tmp | IsNaN_6U_10U_9_nor_3_tmp;
  assign or_967_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | IsNaN_6U_10U_8_land_lpi_1_dfm_4
      | or_tmp_753;
  assign mux_618_nl = MUX_s_1_2_2((or_967_nl), (or_964_nl), or_181_cse);
  assign or_970_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp
      | (~(IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_1_tmp & IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_1_tmp));
  assign or_971_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_12_land_2_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_15_land_2_lpi_1_dfm_4) | IsNaN_6U_10U_10_land_2_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_2_lpi_1_dfm_st;
  assign mux_619_nl = MUX_s_1_2_2((or_971_nl), (or_970_nl), or_181_cse);
  assign or_974_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp
      | (~(IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_2_tmp & IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_2_tmp));
  assign or_975_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_12_land_3_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_15_land_3_lpi_1_dfm_4) | IsNaN_6U_10U_10_land_3_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_3_lpi_1_dfm_st;
  assign mux_620_nl = MUX_s_1_2_2((or_975_nl), (or_974_nl), or_181_cse);
  assign or_978_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp
      | (~(IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_3_tmp & IsNaN_6U_10U_11_IsNaN_6U_10U_11_nor_3_tmp));
  assign or_979_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_12_land_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_15_land_lpi_1_dfm_4) | IsNaN_6U_10U_10_land_lpi_1_dfm_4 |
      IsNaN_6U_10U_14_land_lpi_1_dfm_st;
  assign mux_621_nl = MUX_s_1_2_2((or_979_nl), (or_978_nl), or_181_cse);
  assign mux_623_nl = MUX_s_1_2_2(or_tmp_963, mux_tmp_622, IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp);
  assign nand_73_nl = ~(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_1_tmp & (~ or_tmp_966));
  assign mux_624_nl = MUX_s_1_2_2((nand_73_nl), (mux_623_nl), IsNaN_6U_10U_14_land_2_lpi_1_dfm_st);
  assign mux_625_nl = MUX_s_1_2_2(or_tmp_966, mux_tmp_622, IsNaN_6U_10U_14_land_3_lpi_1_dfm_st);
  assign or_985_nl = (~ IsNaN_6U_10U_14_land_3_lpi_1_dfm_st) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt | (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign mux_626_nl = MUX_s_1_2_2((or_985_nl), (mux_625_nl), IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_2_tmp);
  assign mux_627_nl = MUX_s_1_2_2(or_tmp_966, mux_tmp_622, IsNaN_6U_10U_14_land_lpi_1_dfm_st);
  assign or_986_nl = (~ IsNaN_6U_10U_14_land_lpi_1_dfm_st) | (~ reg_chn_data_out_rsci_ld_core_psct_cse)
      | chn_data_out_rsci_bawt | (~ main_stage_v_2) | m_row0_unequal_tmp_3;
  assign mux_628_nl = MUX_s_1_2_2((or_986_nl), (mux_627_nl), IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_3_tmp);
  assign or_999_nl = (~ IsNaN_6U_10U_12_land_1_lpi_1_dfm_4) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_4
      | (~ reg_chn_data_out_rsci_ld_core_psct_cse) | chn_data_out_rsci_bawt | (~
      main_stage_v_2) | m_row0_unequal_tmp_3;
  assign or_1000_nl = (~ IsNaN_6U_10U_12_land_1_lpi_1_dfm_4) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_4;
  assign mux_639_nl = MUX_s_1_2_2(mux_tmp_622, or_tmp_966, or_1000_nl);
  assign or_998_nl = (~ IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp;
  assign mux_640_nl = MUX_s_1_2_2((mux_639_nl), (or_999_nl), or_998_nl);
  assign or_1003_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp
      | (~(IsNaN_6U_10U_15_IsNaN_6U_10U_15_nor_tmp & IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp));
  assign or_1004_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_12_land_1_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_15_land_1_lpi_1_dfm_4) | IsNaN_6U_10U_10_land_1_lpi_1_dfm_4
      | IsNaN_6U_10U_14_land_1_lpi_1_dfm_st;
  assign mux_641_nl = MUX_s_1_2_2((or_1004_nl), (or_1003_nl), or_181_cse);
  assign or_1006_nl = (cfg_precision!=2'b10) | (~ main_stage_v_1) | (~ IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp)
      | (~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp) | IsNaN_6U_10U_9_IsNaN_6U_10U_9_nor_tmp;
  assign or_1007_nl = (~ main_stage_v_2) | m_row0_unequal_tmp_3 | (~ IsNaN_6U_10U_13_land_1_lpi_1_dfm_4)
      | (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_4) | (~ IsNaN_6U_10U_10_land_1_lpi_1_dfm_4)
      | IsNaN_6U_10U_12_land_1_lpi_1_dfm_4;
  assign mux_642_nl = MUX_s_1_2_2((or_1007_nl), (or_1006_nl), or_181_cse);
  assign mux_643_nl = MUX_s_1_2_2(or_tmp_963, mux_tmp_622, IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp);
  assign nand_77_nl = ~(IsNaN_6U_10U_10_IsNaN_6U_10U_10_nor_tmp & (~ or_tmp_966));
  assign mux_644_nl = MUX_s_1_2_2((nand_77_nl), (mux_643_nl), IsNaN_6U_10U_14_land_1_lpi_1_dfm_st);
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_160_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_sva_1_20_2_1[0])
      & data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_sva_1_20_2_1[0])
      & data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_161_nl = MUX_s_1_2_2((data_truncate_16_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_16_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out = (IntShiftRight_18U_2U_8U_obits_fixed_mux_160_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_161_nl);
  assign z_out = nl_z_out[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_162_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_15_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_1_sva_1_20_2_1[0])
      & data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_15_sva_1_20_2_1[0])
      & data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_163_nl = MUX_s_1_2_2((data_truncate_15_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_1_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_1 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_162_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_163_nl);
  assign z_out_1 = nl_z_out_1[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_164_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_14_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_2_sva_1_20_2_1[0])
      & data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_14_sva_1_20_2_1[0])
      & data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_165_nl = MUX_s_1_2_2((data_truncate_14_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_2_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_2 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_164_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_165_nl);
  assign z_out_2 = nl_z_out_2[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_166_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_13_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_3_sva_1_20_2_1[0])
      & data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_13_sva_1_20_2_1[0])
      & data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_167_nl = MUX_s_1_2_2((data_truncate_13_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_3_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_3 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_166_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_167_nl);
  assign z_out_3 = nl_z_out_3[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_168_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_12_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_4_sva_1_20_2_1[0])
      & data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_12_sva_1_20_2_1[0])
      & data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_169_nl = MUX_s_1_2_2((data_truncate_12_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_4_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_4 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_168_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_169_nl);
  assign z_out_4 = nl_z_out_4[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_170_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_11_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_5_sva_1_20_2_1[0])
      & data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_11_sva_1_20_2_1[0])
      & data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_171_nl = MUX_s_1_2_2((data_truncate_11_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_5_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_5 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_170_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_171_nl);
  assign z_out_5 = nl_z_out_5[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_172_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_10_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_6_sva_1_20_2_1[0])
      & data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_10_sva_1_20_2_1[0])
      & data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_173_nl = MUX_s_1_2_2((data_truncate_10_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_6_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_6 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_172_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_173_nl);
  assign z_out_6 = nl_z_out_6[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_174_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_9_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_7_sva_1_20_2_1[0])
      & data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_9_sva_1_20_2_1[0])
      & data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_175_nl = MUX_s_1_2_2((data_truncate_9_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_7_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_7 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_174_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_175_nl);
  assign z_out_7 = nl_z_out_7[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_176_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_8_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_8_sva_1_20_2_1[0])
      & data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_8_sva_1_20_2_1[0])
      & data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_177_nl = MUX_s_1_2_2((data_truncate_8_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_8_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_8 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_176_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_177_nl);
  assign z_out_8 = nl_z_out_8[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_178_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_7_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_9_sva_1_20_2_1[0])
      & data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_7_sva_1_20_2_1[0])
      & data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_179_nl = MUX_s_1_2_2((data_truncate_7_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_9_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_9 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_178_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_179_nl);
  assign z_out_9 = nl_z_out_9[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_180_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_6_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_10_sva_1_20_2_1[0])
      & data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_6_sva_1_20_2_1[0])
      & data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_181_nl = MUX_s_1_2_2((data_truncate_6_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_10_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_10 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_180_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_181_nl);
  assign z_out_10 = nl_z_out_10[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_182_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_5_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_11_sva_1_20_2_1[0])
      & data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_5_sva_1_20_2_1[0])
      & data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_183_nl = MUX_s_1_2_2((data_truncate_5_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_11_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_11 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_182_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_183_nl);
  assign z_out_11 = nl_z_out_11[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_184_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_4_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_12_sva_1_20_2_1[0])
      & data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_4_sva_1_20_2_1[0])
      & data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_185_nl = MUX_s_1_2_2((data_truncate_4_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_12_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_12 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_184_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_185_nl);
  assign z_out_12 = nl_z_out_12[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_186_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_3_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_13_sva_1_20_2_1[0])
      & data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_3_sva_1_20_2_1[0])
      & data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_187_nl = MUX_s_1_2_2((data_truncate_3_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_13_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_13 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_186_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_187_nl);
  assign z_out_13 = nl_z_out_13[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_188_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_2_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_14_sva_1_20_2_1[0])
      & data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_2_sva_1_20_2_1[0])
      & data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_189_nl = MUX_s_1_2_2((data_truncate_2_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_14_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_14 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_188_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_189_nl);
  assign z_out_14 = nl_z_out_14[17:0];
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_190_nl = MUX_v_18_2_2((IntShiftRight_18U_2U_8U_mbits_fixed_1_sva_1_20_2_1[18:1]),
      (IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_1_20_2_1[18:1]), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_16U_mbits_fixed_15_sva_1_20_2_1[0])
      & data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_or_itm_2;
  assign data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl = (IntShiftRight_18U_2U_8U_mbits_fixed_1_sva_1_20_2_1[0])
      & data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_or_itm_2;
  assign IntShiftRight_18U_2U_8U_obits_fixed_mux_191_nl = MUX_s_1_2_2((data_truncate_1_IntShiftRight_18U_2U_8U_obits_fixed_and_2_nl),
      (data_truncate_15_IntShiftRight_18U_2U_16U_obits_fixed_and_2_nl), IntShiftRight_18U_2U_16U_obits_fixed_and_111_cse);
  assign nl_z_out_15 = (IntShiftRight_18U_2U_8U_obits_fixed_mux_190_nl) + conv_u2u_1_18(IntShiftRight_18U_2U_8U_obits_fixed_mux_191_nl);
  assign z_out_15 = nl_z_out_15[17:0];

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction


  function [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    result = result | ( input_4 & {6{sel[4]}});
    result = result | ( input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction


  function [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function [23:0] readslicef_25_24_1;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_25_24_1 = tmp[23:0];
  end
  endfunction


  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function  [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function  [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function  [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function  [9:0] conv_u2u_1_10 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [10:0] conv_u2u_1_11 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction


  function  [17:0] conv_u2u_1_18 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_18 = {{17{1'b0}}, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function  [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function  [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function  [23:0] conv_u2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_u2u_23_24 = {1'b0, vector};
  end
  endfunction


  function  [24:0] conv_u2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_u2u_24_25 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    NV_NVDLA_CSC_pra_cell
// ------------------------------------------------------------------


module NV_NVDLA_CSC_pra_cell (
  nvdla_core_clk, nvdla_core_rstn, chn_data_in_rsc_z, chn_data_in_rsc_vz, chn_data_in_rsc_lz,
      cfg_precision, cfg_truncate_rsc_z, chn_data_out_rsc_z, chn_data_out_rsc_vz,
      chn_data_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [255:0] chn_data_in_rsc_z;
  input chn_data_in_rsc_vz;
  output chn_data_in_rsc_lz;
  input [1:0] cfg_precision;
  input [1:0] cfg_truncate_rsc_z;
  output [255:0] chn_data_out_rsc_z;
  input chn_data_out_rsc_vz;
  output chn_data_out_rsc_lz;


  // Interconnect Declarations
  wire chn_data_in_rsci_oswt;
  wire chn_data_in_rsci_oswt_unreg;
  wire chn_data_out_rsci_oswt;
  wire chn_data_out_rsci_oswt_unreg;


  // Interconnect Declarations for Component Instantiations 
  CSC_chn_data_in_rsci_unreg chn_data_in_rsci_unreg_inst (
      .in_0(chn_data_in_rsci_oswt_unreg),
      .outsig(chn_data_in_rsci_oswt)
    );
  CSC_chn_data_out_rsci_unreg chn_data_out_rsci_unreg_inst (
      .in_0(chn_data_out_rsci_oswt_unreg),
      .outsig(chn_data_out_rsci_oswt)
    );
  NV_NVDLA_CSC_pra_cell_core NV_NVDLA_CSC_pra_cell_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_data_in_rsc_z(chn_data_in_rsc_z),
      .chn_data_in_rsc_vz(chn_data_in_rsc_vz),
      .chn_data_in_rsc_lz(chn_data_in_rsc_lz),
      .cfg_precision(cfg_precision),
      .cfg_truncate_rsc_z(cfg_truncate_rsc_z),
      .chn_data_out_rsc_z(chn_data_out_rsc_z),
      .chn_data_out_rsc_vz(chn_data_out_rsc_vz),
      .chn_data_out_rsc_lz(chn_data_out_rsc_lz),
      .chn_data_in_rsci_oswt(chn_data_in_rsci_oswt),
      .chn_data_in_rsci_oswt_unreg(chn_data_in_rsci_oswt_unreg),
      .chn_data_out_rsci_oswt(chn_data_out_rsci_oswt),
      .chn_data_out_rsci_oswt_unreg(chn_data_out_rsci_oswt_unreg)
    );
endmodule



