// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_NVDLA_CMAC_CORE_active.v

module NV_NVDLA_CMAC_CORE_active (
   nvdla_core_clk
  ,nvdla_core_rstn
  ,cfg_is_fp16
  ,cfg_is_int16
  ,cfg_is_int8
  ,cfg_reg_en
  ,in_dat_data0
  ,in_dat_data1
  ,in_dat_data10
  ,in_dat_data100
  ,in_dat_data101
  ,in_dat_data102
  ,in_dat_data103
  ,in_dat_data104
  ,in_dat_data105
  ,in_dat_data106
  ,in_dat_data107
  ,in_dat_data108
  ,in_dat_data109
  ,in_dat_data11
  ,in_dat_data110
  ,in_dat_data111
  ,in_dat_data112
  ,in_dat_data113
  ,in_dat_data114
  ,in_dat_data115
  ,in_dat_data116
  ,in_dat_data117
  ,in_dat_data118
  ,in_dat_data119
  ,in_dat_data12
  ,in_dat_data120
  ,in_dat_data121
  ,in_dat_data122
  ,in_dat_data123
  ,in_dat_data124
  ,in_dat_data125
  ,in_dat_data126
  ,in_dat_data127
  ,in_dat_data13
  ,in_dat_data14
  ,in_dat_data15
  ,in_dat_data16
  ,in_dat_data17
  ,in_dat_data18
  ,in_dat_data19
  ,in_dat_data2
  ,in_dat_data20
  ,in_dat_data21
  ,in_dat_data22
  ,in_dat_data23
  ,in_dat_data24
  ,in_dat_data25
  ,in_dat_data26
  ,in_dat_data27
  ,in_dat_data28
  ,in_dat_data29
  ,in_dat_data3
  ,in_dat_data30
  ,in_dat_data31
  ,in_dat_data32
  ,in_dat_data33
  ,in_dat_data34
  ,in_dat_data35
  ,in_dat_data36
  ,in_dat_data37
  ,in_dat_data38
  ,in_dat_data39
  ,in_dat_data4
  ,in_dat_data40
  ,in_dat_data41
  ,in_dat_data42
  ,in_dat_data43
  ,in_dat_data44
  ,in_dat_data45
  ,in_dat_data46
  ,in_dat_data47
  ,in_dat_data48
  ,in_dat_data49
  ,in_dat_data5
  ,in_dat_data50
  ,in_dat_data51
  ,in_dat_data52
  ,in_dat_data53
  ,in_dat_data54
  ,in_dat_data55
  ,in_dat_data56
  ,in_dat_data57
  ,in_dat_data58
  ,in_dat_data59
  ,in_dat_data6
  ,in_dat_data60
  ,in_dat_data61
  ,in_dat_data62
  ,in_dat_data63
  ,in_dat_data64
  ,in_dat_data65
  ,in_dat_data66
  ,in_dat_data67
  ,in_dat_data68
  ,in_dat_data69
  ,in_dat_data7
  ,in_dat_data70
  ,in_dat_data71
  ,in_dat_data72
  ,in_dat_data73
  ,in_dat_data74
  ,in_dat_data75
  ,in_dat_data76
  ,in_dat_data77
  ,in_dat_data78
  ,in_dat_data79
  ,in_dat_data8
  ,in_dat_data80
  ,in_dat_data81
  ,in_dat_data82
  ,in_dat_data83
  ,in_dat_data84
  ,in_dat_data85
  ,in_dat_data86
  ,in_dat_data87
  ,in_dat_data88
  ,in_dat_data89
  ,in_dat_data9
  ,in_dat_data90
  ,in_dat_data91
  ,in_dat_data92
  ,in_dat_data93
  ,in_dat_data94
  ,in_dat_data95
  ,in_dat_data96
  ,in_dat_data97
  ,in_dat_data98
  ,in_dat_data99
  ,in_dat_mask
  ,in_dat_pvld
  ,in_dat_stripe_end
  ,in_dat_stripe_st
  ,in_wt_data0
  ,in_wt_data1
  ,in_wt_data10
  ,in_wt_data100
  ,in_wt_data101
  ,in_wt_data102
  ,in_wt_data103
  ,in_wt_data104
  ,in_wt_data105
  ,in_wt_data106
  ,in_wt_data107
  ,in_wt_data108
  ,in_wt_data109
  ,in_wt_data11
  ,in_wt_data110
  ,in_wt_data111
  ,in_wt_data112
  ,in_wt_data113
  ,in_wt_data114
  ,in_wt_data115
  ,in_wt_data116
  ,in_wt_data117
  ,in_wt_data118
  ,in_wt_data119
  ,in_wt_data12
  ,in_wt_data120
  ,in_wt_data121
  ,in_wt_data122
  ,in_wt_data123
  ,in_wt_data124
  ,in_wt_data125
  ,in_wt_data126
  ,in_wt_data127
  ,in_wt_data13
  ,in_wt_data14
  ,in_wt_data15
  ,in_wt_data16
  ,in_wt_data17
  ,in_wt_data18
  ,in_wt_data19
  ,in_wt_data2
  ,in_wt_data20
  ,in_wt_data21
  ,in_wt_data22
  ,in_wt_data23
  ,in_wt_data24
  ,in_wt_data25
  ,in_wt_data26
  ,in_wt_data27
  ,in_wt_data28
  ,in_wt_data29
  ,in_wt_data3
  ,in_wt_data30
  ,in_wt_data31
  ,in_wt_data32
  ,in_wt_data33
  ,in_wt_data34
  ,in_wt_data35
  ,in_wt_data36
  ,in_wt_data37
  ,in_wt_data38
  ,in_wt_data39
  ,in_wt_data4
  ,in_wt_data40
  ,in_wt_data41
  ,in_wt_data42
  ,in_wt_data43
  ,in_wt_data44
  ,in_wt_data45
  ,in_wt_data46
  ,in_wt_data47
  ,in_wt_data48
  ,in_wt_data49
  ,in_wt_data5
  ,in_wt_data50
  ,in_wt_data51
  ,in_wt_data52
  ,in_wt_data53
  ,in_wt_data54
  ,in_wt_data55
  ,in_wt_data56
  ,in_wt_data57
  ,in_wt_data58
  ,in_wt_data59
  ,in_wt_data6
  ,in_wt_data60
  ,in_wt_data61
  ,in_wt_data62
  ,in_wt_data63
  ,in_wt_data64
  ,in_wt_data65
  ,in_wt_data66
  ,in_wt_data67
  ,in_wt_data68
  ,in_wt_data69
  ,in_wt_data7
  ,in_wt_data70
  ,in_wt_data71
  ,in_wt_data72
  ,in_wt_data73
  ,in_wt_data74
  ,in_wt_data75
  ,in_wt_data76
  ,in_wt_data77
  ,in_wt_data78
  ,in_wt_data79
  ,in_wt_data8
  ,in_wt_data80
  ,in_wt_data81
  ,in_wt_data82
  ,in_wt_data83
  ,in_wt_data84
  ,in_wt_data85
  ,in_wt_data86
  ,in_wt_data87
  ,in_wt_data88
  ,in_wt_data89
  ,in_wt_data9
  ,in_wt_data90
  ,in_wt_data91
  ,in_wt_data92
  ,in_wt_data93
  ,in_wt_data94
  ,in_wt_data95
  ,in_wt_data96
  ,in_wt_data97
  ,in_wt_data98
  ,in_wt_data99
  ,in_wt_mask
  ,in_wt_pvld
  ,in_wt_sel
  ,dat0_actv_data
  ,dat0_actv_nan
  ,dat0_actv_nz
  ,dat0_actv_pvld
  ,dat0_pre_exp
  ,dat0_pre_mask
  ,dat0_pre_pvld
  ,dat0_pre_stripe_end
  ,dat0_pre_stripe_st
  ,dat1_actv_data
  ,dat1_actv_nan
  ,dat1_actv_nz
  ,dat1_actv_pvld
  ,dat1_pre_exp
  ,dat1_pre_mask
  ,dat1_pre_pvld
  ,dat1_pre_stripe_end
  ,dat1_pre_stripe_st
  ,dat2_actv_data
  ,dat2_actv_nan
  ,dat2_actv_nz
  ,dat2_actv_pvld
  ,dat2_pre_exp
  ,dat2_pre_mask
  ,dat2_pre_pvld
  ,dat2_pre_stripe_end
  ,dat2_pre_stripe_st
  ,dat3_actv_data
  ,dat3_actv_nan
  ,dat3_actv_nz
  ,dat3_actv_pvld
  ,dat3_pre_exp
  ,dat3_pre_mask
  ,dat3_pre_pvld
  ,dat3_pre_stripe_end
  ,dat3_pre_stripe_st
  ,dat4_actv_data
  ,dat4_actv_nan
  ,dat4_actv_nz
  ,dat4_actv_pvld
  ,dat4_pre_exp
  ,dat4_pre_mask
  ,dat4_pre_pvld
  ,dat4_pre_stripe_end
  ,dat4_pre_stripe_st
  ,dat5_actv_data
  ,dat5_actv_nan
  ,dat5_actv_nz
  ,dat5_actv_pvld
  ,dat5_pre_exp
  ,dat5_pre_mask
  ,dat5_pre_pvld
  ,dat5_pre_stripe_end
  ,dat5_pre_stripe_st
  ,dat6_actv_data
  ,dat6_actv_nan
  ,dat6_actv_nz
  ,dat6_actv_pvld
  ,dat6_pre_exp
  ,dat6_pre_mask
  ,dat6_pre_pvld
  ,dat6_pre_stripe_end
  ,dat6_pre_stripe_st
  ,dat7_actv_data
  ,dat7_actv_nan
  ,dat7_actv_nz
  ,dat7_actv_pvld
  ,dat7_pre_exp
  ,dat7_pre_mask
  ,dat7_pre_pvld
  ,dat7_pre_stripe_end
  ,dat7_pre_stripe_st
  ,wt0_actv_data
  ,wt0_actv_nan
  ,wt0_actv_nz
  ,wt0_actv_pvld
  ,wt0_sd_exp
  ,wt0_sd_mask
  ,wt0_sd_pvld
  ,wt1_actv_data
  ,wt1_actv_nan
  ,wt1_actv_nz
  ,wt1_actv_pvld
  ,wt1_sd_exp
  ,wt1_sd_mask
  ,wt1_sd_pvld
  ,wt2_actv_data
  ,wt2_actv_nan
  ,wt2_actv_nz
  ,wt2_actv_pvld
  ,wt2_sd_exp
  ,wt2_sd_mask
  ,wt2_sd_pvld
  ,wt3_actv_data
  ,wt3_actv_nan
  ,wt3_actv_nz
  ,wt3_actv_pvld
  ,wt3_sd_exp
  ,wt3_sd_mask
  ,wt3_sd_pvld
  ,wt4_actv_data
  ,wt4_actv_nan
  ,wt4_actv_nz
  ,wt4_actv_pvld
  ,wt4_sd_exp
  ,wt4_sd_mask
  ,wt4_sd_pvld
  ,wt5_actv_data
  ,wt5_actv_nan
  ,wt5_actv_nz
  ,wt5_actv_pvld
  ,wt5_sd_exp
  ,wt5_sd_mask
  ,wt5_sd_pvld
  ,wt6_actv_data
  ,wt6_actv_nan
  ,wt6_actv_nz
  ,wt6_actv_pvld
  ,wt6_sd_exp
  ,wt6_sd_mask
  ,wt6_sd_pvld
  ,wt7_actv_data
  ,wt7_actv_nan
  ,wt7_actv_nz
  ,wt7_actv_pvld
  ,wt7_sd_exp
  ,wt7_sd_mask
  ,wt7_sd_pvld
  );

input           nvdla_core_clk;
input           nvdla_core_rstn;
input           cfg_is_fp16;
input           cfg_is_int16;
input           cfg_is_int8;
input           cfg_reg_en;
input     [7:0] in_dat_data0;
input     [7:0] in_dat_data1;
input     [7:0] in_dat_data10;
input     [7:0] in_dat_data100;
input     [7:0] in_dat_data101;
input     [7:0] in_dat_data102;
input     [7:0] in_dat_data103;
input     [7:0] in_dat_data104;
input     [7:0] in_dat_data105;
input     [7:0] in_dat_data106;
input     [7:0] in_dat_data107;
input     [7:0] in_dat_data108;
input     [7:0] in_dat_data109;
input     [7:0] in_dat_data11;
input     [7:0] in_dat_data110;
input     [7:0] in_dat_data111;
input     [7:0] in_dat_data112;
input     [7:0] in_dat_data113;
input     [7:0] in_dat_data114;
input     [7:0] in_dat_data115;
input     [7:0] in_dat_data116;
input     [7:0] in_dat_data117;
input     [7:0] in_dat_data118;
input     [7:0] in_dat_data119;
input     [7:0] in_dat_data12;
input     [7:0] in_dat_data120;
input     [7:0] in_dat_data121;
input     [7:0] in_dat_data122;
input     [7:0] in_dat_data123;
input     [7:0] in_dat_data124;
input     [7:0] in_dat_data125;
input     [7:0] in_dat_data126;
input     [7:0] in_dat_data127;
input     [7:0] in_dat_data13;
input     [7:0] in_dat_data14;
input     [7:0] in_dat_data15;
input     [7:0] in_dat_data16;
input     [7:0] in_dat_data17;
input     [7:0] in_dat_data18;
input     [7:0] in_dat_data19;
input     [7:0] in_dat_data2;
input     [7:0] in_dat_data20;
input     [7:0] in_dat_data21;
input     [7:0] in_dat_data22;
input     [7:0] in_dat_data23;
input     [7:0] in_dat_data24;
input     [7:0] in_dat_data25;
input     [7:0] in_dat_data26;
input     [7:0] in_dat_data27;
input     [7:0] in_dat_data28;
input     [7:0] in_dat_data29;
input     [7:0] in_dat_data3;
input     [7:0] in_dat_data30;
input     [7:0] in_dat_data31;
input     [7:0] in_dat_data32;
input     [7:0] in_dat_data33;
input     [7:0] in_dat_data34;
input     [7:0] in_dat_data35;
input     [7:0] in_dat_data36;
input     [7:0] in_dat_data37;
input     [7:0] in_dat_data38;
input     [7:0] in_dat_data39;
input     [7:0] in_dat_data4;
input     [7:0] in_dat_data40;
input     [7:0] in_dat_data41;
input     [7:0] in_dat_data42;
input     [7:0] in_dat_data43;
input     [7:0] in_dat_data44;
input     [7:0] in_dat_data45;
input     [7:0] in_dat_data46;
input     [7:0] in_dat_data47;
input     [7:0] in_dat_data48;
input     [7:0] in_dat_data49;
input     [7:0] in_dat_data5;
input     [7:0] in_dat_data50;
input     [7:0] in_dat_data51;
input     [7:0] in_dat_data52;
input     [7:0] in_dat_data53;
input     [7:0] in_dat_data54;
input     [7:0] in_dat_data55;
input     [7:0] in_dat_data56;
input     [7:0] in_dat_data57;
input     [7:0] in_dat_data58;
input     [7:0] in_dat_data59;
input     [7:0] in_dat_data6;
input     [7:0] in_dat_data60;
input     [7:0] in_dat_data61;
input     [7:0] in_dat_data62;
input     [7:0] in_dat_data63;
input     [7:0] in_dat_data64;
input     [7:0] in_dat_data65;
input     [7:0] in_dat_data66;
input     [7:0] in_dat_data67;
input     [7:0] in_dat_data68;
input     [7:0] in_dat_data69;
input     [7:0] in_dat_data7;
input     [7:0] in_dat_data70;
input     [7:0] in_dat_data71;
input     [7:0] in_dat_data72;
input     [7:0] in_dat_data73;
input     [7:0] in_dat_data74;
input     [7:0] in_dat_data75;
input     [7:0] in_dat_data76;
input     [7:0] in_dat_data77;
input     [7:0] in_dat_data78;
input     [7:0] in_dat_data79;
input     [7:0] in_dat_data8;
input     [7:0] in_dat_data80;
input     [7:0] in_dat_data81;
input     [7:0] in_dat_data82;
input     [7:0] in_dat_data83;
input     [7:0] in_dat_data84;
input     [7:0] in_dat_data85;
input     [7:0] in_dat_data86;
input     [7:0] in_dat_data87;
input     [7:0] in_dat_data88;
input     [7:0] in_dat_data89;
input     [7:0] in_dat_data9;
input     [7:0] in_dat_data90;
input     [7:0] in_dat_data91;
input     [7:0] in_dat_data92;
input     [7:0] in_dat_data93;
input     [7:0] in_dat_data94;
input     [7:0] in_dat_data95;
input     [7:0] in_dat_data96;
input     [7:0] in_dat_data97;
input     [7:0] in_dat_data98;
input     [7:0] in_dat_data99;
input   [127:0] in_dat_mask;
input           in_dat_pvld;
input           in_dat_stripe_end;
input           in_dat_stripe_st;
input     [7:0] in_wt_data0;
input     [7:0] in_wt_data1;
input     [7:0] in_wt_data10;
input     [7:0] in_wt_data100;
input     [7:0] in_wt_data101;
input     [7:0] in_wt_data102;
input     [7:0] in_wt_data103;
input     [7:0] in_wt_data104;
input     [7:0] in_wt_data105;
input     [7:0] in_wt_data106;
input     [7:0] in_wt_data107;
input     [7:0] in_wt_data108;
input     [7:0] in_wt_data109;
input     [7:0] in_wt_data11;
input     [7:0] in_wt_data110;
input     [7:0] in_wt_data111;
input     [7:0] in_wt_data112;
input     [7:0] in_wt_data113;
input     [7:0] in_wt_data114;
input     [7:0] in_wt_data115;
input     [7:0] in_wt_data116;
input     [7:0] in_wt_data117;
input     [7:0] in_wt_data118;
input     [7:0] in_wt_data119;
input     [7:0] in_wt_data12;
input     [7:0] in_wt_data120;
input     [7:0] in_wt_data121;
input     [7:0] in_wt_data122;
input     [7:0] in_wt_data123;
input     [7:0] in_wt_data124;
input     [7:0] in_wt_data125;
input     [7:0] in_wt_data126;
input     [7:0] in_wt_data127;
input     [7:0] in_wt_data13;
input     [7:0] in_wt_data14;
input     [7:0] in_wt_data15;
input     [7:0] in_wt_data16;
input     [7:0] in_wt_data17;
input     [7:0] in_wt_data18;
input     [7:0] in_wt_data19;
input     [7:0] in_wt_data2;
input     [7:0] in_wt_data20;
input     [7:0] in_wt_data21;
input     [7:0] in_wt_data22;
input     [7:0] in_wt_data23;
input     [7:0] in_wt_data24;
input     [7:0] in_wt_data25;
input     [7:0] in_wt_data26;
input     [7:0] in_wt_data27;
input     [7:0] in_wt_data28;
input     [7:0] in_wt_data29;
input     [7:0] in_wt_data3;
input     [7:0] in_wt_data30;
input     [7:0] in_wt_data31;
input     [7:0] in_wt_data32;
input     [7:0] in_wt_data33;
input     [7:0] in_wt_data34;
input     [7:0] in_wt_data35;
input     [7:0] in_wt_data36;
input     [7:0] in_wt_data37;
input     [7:0] in_wt_data38;
input     [7:0] in_wt_data39;
input     [7:0] in_wt_data4;
input     [7:0] in_wt_data40;
input     [7:0] in_wt_data41;
input     [7:0] in_wt_data42;
input     [7:0] in_wt_data43;
input     [7:0] in_wt_data44;
input     [7:0] in_wt_data45;
input     [7:0] in_wt_data46;
input     [7:0] in_wt_data47;
input     [7:0] in_wt_data48;
input     [7:0] in_wt_data49;
input     [7:0] in_wt_data5;
input     [7:0] in_wt_data50;
input     [7:0] in_wt_data51;
input     [7:0] in_wt_data52;
input     [7:0] in_wt_data53;
input     [7:0] in_wt_data54;
input     [7:0] in_wt_data55;
input     [7:0] in_wt_data56;
input     [7:0] in_wt_data57;
input     [7:0] in_wt_data58;
input     [7:0] in_wt_data59;
input     [7:0] in_wt_data6;
input     [7:0] in_wt_data60;
input     [7:0] in_wt_data61;
input     [7:0] in_wt_data62;
input     [7:0] in_wt_data63;
input     [7:0] in_wt_data64;
input     [7:0] in_wt_data65;
input     [7:0] in_wt_data66;
input     [7:0] in_wt_data67;
input     [7:0] in_wt_data68;
input     [7:0] in_wt_data69;
input     [7:0] in_wt_data7;
input     [7:0] in_wt_data70;
input     [7:0] in_wt_data71;
input     [7:0] in_wt_data72;
input     [7:0] in_wt_data73;
input     [7:0] in_wt_data74;
input     [7:0] in_wt_data75;
input     [7:0] in_wt_data76;
input     [7:0] in_wt_data77;
input     [7:0] in_wt_data78;
input     [7:0] in_wt_data79;
input     [7:0] in_wt_data8;
input     [7:0] in_wt_data80;
input     [7:0] in_wt_data81;
input     [7:0] in_wt_data82;
input     [7:0] in_wt_data83;
input     [7:0] in_wt_data84;
input     [7:0] in_wt_data85;
input     [7:0] in_wt_data86;
input     [7:0] in_wt_data87;
input     [7:0] in_wt_data88;
input     [7:0] in_wt_data89;
input     [7:0] in_wt_data9;
input     [7:0] in_wt_data90;
input     [7:0] in_wt_data91;
input     [7:0] in_wt_data92;
input     [7:0] in_wt_data93;
input     [7:0] in_wt_data94;
input     [7:0] in_wt_data95;
input     [7:0] in_wt_data96;
input     [7:0] in_wt_data97;
input     [7:0] in_wt_data98;
input     [7:0] in_wt_data99;
input   [127:0] in_wt_mask;
input           in_wt_pvld;
input     [7:0] in_wt_sel;
output [1023:0] dat0_actv_data;
output   [63:0] dat0_actv_nan;
output  [127:0] dat0_actv_nz;
output  [103:0] dat0_actv_pvld;
output  [191:0] dat0_pre_exp;
output   [63:0] dat0_pre_mask;
output          dat0_pre_pvld;
output          dat0_pre_stripe_end;
output          dat0_pre_stripe_st;
output [1023:0] dat1_actv_data;
output   [63:0] dat1_actv_nan;
output  [127:0] dat1_actv_nz;
output  [103:0] dat1_actv_pvld;
output  [191:0] dat1_pre_exp;
output   [63:0] dat1_pre_mask;
output          dat1_pre_pvld;
output          dat1_pre_stripe_end;
output          dat1_pre_stripe_st;
output [1023:0] dat2_actv_data;
output   [63:0] dat2_actv_nan;
output  [127:0] dat2_actv_nz;
output  [103:0] dat2_actv_pvld;
output  [191:0] dat2_pre_exp;
output   [63:0] dat2_pre_mask;
output          dat2_pre_pvld;
output          dat2_pre_stripe_end;
output          dat2_pre_stripe_st;
output [1023:0] dat3_actv_data;
output   [63:0] dat3_actv_nan;
output  [127:0] dat3_actv_nz;
output  [103:0] dat3_actv_pvld;
output  [191:0] dat3_pre_exp;
output   [63:0] dat3_pre_mask;
output          dat3_pre_pvld;
output          dat3_pre_stripe_end;
output          dat3_pre_stripe_st;
output [1023:0] dat4_actv_data;
output   [63:0] dat4_actv_nan;
output  [127:0] dat4_actv_nz;
output  [103:0] dat4_actv_pvld;
output  [191:0] dat4_pre_exp;
output   [63:0] dat4_pre_mask;
output          dat4_pre_pvld;
output          dat4_pre_stripe_end;
output          dat4_pre_stripe_st;
output [1023:0] dat5_actv_data;
output   [63:0] dat5_actv_nan;
output  [127:0] dat5_actv_nz;
output  [103:0] dat5_actv_pvld;
output  [191:0] dat5_pre_exp;
output   [63:0] dat5_pre_mask;
output          dat5_pre_pvld;
output          dat5_pre_stripe_end;
output          dat5_pre_stripe_st;
output [1023:0] dat6_actv_data;
output   [63:0] dat6_actv_nan;
output  [127:0] dat6_actv_nz;
output  [103:0] dat6_actv_pvld;
output  [191:0] dat6_pre_exp;
output   [63:0] dat6_pre_mask;
output          dat6_pre_pvld;
output          dat6_pre_stripe_end;
output          dat6_pre_stripe_st;
output [1023:0] dat7_actv_data;
output   [63:0] dat7_actv_nan;
output  [127:0] dat7_actv_nz;
output  [103:0] dat7_actv_pvld;
output  [191:0] dat7_pre_exp;
output   [63:0] dat7_pre_mask;
output          dat7_pre_pvld;
output          dat7_pre_stripe_end;
output          dat7_pre_stripe_st;
output [1023:0] wt0_actv_data;
output   [63:0] wt0_actv_nan;
output  [127:0] wt0_actv_nz;
output  [103:0] wt0_actv_pvld;
output  [191:0] wt0_sd_exp;
output   [63:0] wt0_sd_mask;
output          wt0_sd_pvld;
output [1023:0] wt1_actv_data;
output   [63:0] wt1_actv_nan;
output  [127:0] wt1_actv_nz;
output  [103:0] wt1_actv_pvld;
output  [191:0] wt1_sd_exp;
output   [63:0] wt1_sd_mask;
output          wt1_sd_pvld;
output [1023:0] wt2_actv_data;
output   [63:0] wt2_actv_nan;
output  [127:0] wt2_actv_nz;
output  [103:0] wt2_actv_pvld;
output  [191:0] wt2_sd_exp;
output   [63:0] wt2_sd_mask;
output          wt2_sd_pvld;
output [1023:0] wt3_actv_data;
output   [63:0] wt3_actv_nan;
output  [127:0] wt3_actv_nz;
output  [103:0] wt3_actv_pvld;
output  [191:0] wt3_sd_exp;
output   [63:0] wt3_sd_mask;
output          wt3_sd_pvld;
output [1023:0] wt4_actv_data;
output   [63:0] wt4_actv_nan;
output  [127:0] wt4_actv_nz;
output  [103:0] wt4_actv_pvld;
output  [191:0] wt4_sd_exp;
output   [63:0] wt4_sd_mask;
output          wt4_sd_pvld;
output [1023:0] wt5_actv_data;
output   [63:0] wt5_actv_nan;
output  [127:0] wt5_actv_nz;
output  [103:0] wt5_actv_pvld;
output  [191:0] wt5_sd_exp;
output   [63:0] wt5_sd_mask;
output          wt5_sd_pvld;
output [1023:0] wt6_actv_data;
output   [63:0] wt6_actv_nan;
output  [127:0] wt6_actv_nz;
output  [103:0] wt6_actv_pvld;
output  [191:0] wt6_sd_exp;
output   [63:0] wt6_sd_mask;
output          wt6_sd_pvld;
output [1023:0] wt7_actv_data;
output   [63:0] wt7_actv_nan;
output  [127:0] wt7_actv_nz;
output  [103:0] wt7_actv_pvld;
output  [191:0] wt7_sd_exp;
output   [63:0] wt7_sd_mask;
output          wt7_sd_pvld;
reg      [97:0] cfg_is_fp16_d1;
reg      [63:0] cfg_is_int16_d1;
reg      [64:0] cfg_is_int8_d1;
reg    [1023:0] dat0_actv_data;
reg      [63:0] dat0_actv_nan;
reg     [127:0] dat0_actv_nz;
reg     [103:0] dat0_actv_pvld;
reg     [191:0] dat0_pre_exp;
reg      [63:0] dat0_pre_mask;
reg             dat0_pre_pvld;
reg             dat0_pre_stripe_end;
reg             dat0_pre_stripe_st;
reg    [1023:0] dat1_actv_data;
reg      [63:0] dat1_actv_nan;
reg     [127:0] dat1_actv_nz;
reg     [103:0] dat1_actv_pvld;
reg     [191:0] dat1_pre_exp;
reg      [63:0] dat1_pre_mask;
reg             dat1_pre_pvld;
reg             dat1_pre_stripe_end;
reg             dat1_pre_stripe_st;
reg    [1023:0] dat2_actv_data;
reg      [63:0] dat2_actv_nan;
reg     [127:0] dat2_actv_nz;
reg     [103:0] dat2_actv_pvld;
reg     [191:0] dat2_pre_exp;
reg      [63:0] dat2_pre_mask;
reg             dat2_pre_pvld;
reg             dat2_pre_stripe_end;
reg             dat2_pre_stripe_st;
reg    [1023:0] dat3_actv_data;
reg      [63:0] dat3_actv_nan;
reg     [127:0] dat3_actv_nz;
reg     [103:0] dat3_actv_pvld;
reg     [191:0] dat3_pre_exp;
reg      [63:0] dat3_pre_mask;
reg             dat3_pre_pvld;
reg             dat3_pre_stripe_end;
reg             dat3_pre_stripe_st;
reg    [1023:0] dat4_actv_data;
reg      [63:0] dat4_actv_nan;
reg     [127:0] dat4_actv_nz;
reg     [103:0] dat4_actv_pvld;
reg     [191:0] dat4_pre_exp;
reg      [63:0] dat4_pre_mask;
reg             dat4_pre_pvld;
reg             dat4_pre_stripe_end;
reg             dat4_pre_stripe_st;
reg    [1023:0] dat5_actv_data;
reg      [63:0] dat5_actv_nan;
reg     [127:0] dat5_actv_nz;
reg     [103:0] dat5_actv_pvld;
reg     [191:0] dat5_pre_exp;
reg      [63:0] dat5_pre_mask;
reg             dat5_pre_pvld;
reg             dat5_pre_stripe_end;
reg             dat5_pre_stripe_st;
reg    [1023:0] dat6_actv_data;
reg      [63:0] dat6_actv_nan;
reg     [127:0] dat6_actv_nz;
reg     [103:0] dat6_actv_pvld;
reg     [191:0] dat6_pre_exp;
reg      [63:0] dat6_pre_mask;
reg             dat6_pre_pvld;
reg             dat6_pre_stripe_end;
reg             dat6_pre_stripe_st;
reg    [1023:0] dat7_actv_data;
reg      [63:0] dat7_actv_nan;
reg     [127:0] dat7_actv_nz;
reg     [103:0] dat7_actv_pvld;
reg     [191:0] dat7_pre_exp;
reg      [63:0] dat7_pre_mask;
reg             dat7_pre_pvld;
reg             dat7_pre_stripe_end;
reg             dat7_pre_stripe_st;
reg    [1023:0] dat_actv_data_reg0;
reg    [1023:0] dat_actv_data_reg1;
reg    [1023:0] dat_actv_data_reg2;
reg    [1023:0] dat_actv_data_reg3;
reg    [1023:0] dat_actv_data_reg4;
reg    [1023:0] dat_actv_data_reg5;
reg    [1023:0] dat_actv_data_reg6;
reg    [1023:0] dat_actv_data_reg7;
reg      [63:0] dat_actv_nan_reg0;
reg      [63:0] dat_actv_nan_reg1;
reg      [63:0] dat_actv_nan_reg2;
reg      [63:0] dat_actv_nan_reg3;
reg      [63:0] dat_actv_nan_reg4;
reg      [63:0] dat_actv_nan_reg5;
reg      [63:0] dat_actv_nan_reg6;
reg      [63:0] dat_actv_nan_reg7;
reg     [127:0] dat_actv_nz_reg0;
reg     [127:0] dat_actv_nz_reg1;
reg     [127:0] dat_actv_nz_reg2;
reg     [127:0] dat_actv_nz_reg3;
reg     [127:0] dat_actv_nz_reg4;
reg     [127:0] dat_actv_nz_reg5;
reg     [127:0] dat_actv_nz_reg6;
reg     [127:0] dat_actv_nz_reg7;
reg     [103:0] dat_actv_pvld_reg0;
reg     [103:0] dat_actv_pvld_reg1;
reg     [103:0] dat_actv_pvld_reg2;
reg     [103:0] dat_actv_pvld_reg3;
reg     [103:0] dat_actv_pvld_reg4;
reg     [103:0] dat_actv_pvld_reg5;
reg     [103:0] dat_actv_pvld_reg6;
reg     [103:0] dat_actv_pvld_reg7;
reg             dat_actv_stripe_end;
reg             dat_has_nan;
reg    [1023:0] dat_pre_data;
reg    [1023:0] dat_pre_data_w;
reg     [191:0] dat_pre_exp_reg0;
reg     [191:0] dat_pre_exp_reg1;
reg     [191:0] dat_pre_exp_reg2;
reg     [191:0] dat_pre_exp_reg3;
reg     [191:0] dat_pre_exp_reg4;
reg     [191:0] dat_pre_exp_reg5;
reg     [191:0] dat_pre_exp_reg6;
reg     [191:0] dat_pre_exp_reg7;
reg     [191:0] dat_pre_exp_w;
reg      [63:0] dat_pre_mask0;
reg      [63:0] dat_pre_mask1;
reg      [63:0] dat_pre_mask2;
reg      [63:0] dat_pre_mask3;
reg      [63:0] dat_pre_mask4;
reg      [63:0] dat_pre_mask5;
reg      [63:0] dat_pre_mask6;
reg      [63:0] dat_pre_mask7;
reg      [63:0] dat_pre_mask_w;
reg      [63:0] dat_pre_nan;
reg     [127:0] dat_pre_nz;
reg     [127:0] dat_pre_nz_w;
reg      [15:0] dat_pre_pvld;
reg       [8:0] dat_pre_stripe_end;
reg      [15:0] dat_pre_stripe_st;
reg    [1023:0] in_dat_data_fp16;
reg      [15:0] in_dat_data_fp16_0;
reg      [15:0] in_dat_data_fp16_1;
reg      [15:0] in_dat_data_fp16_10;
reg      [15:0] in_dat_data_fp16_11;
reg      [15:0] in_dat_data_fp16_12;
reg      [15:0] in_dat_data_fp16_13;
reg      [15:0] in_dat_data_fp16_14;
reg      [15:0] in_dat_data_fp16_15;
reg      [15:0] in_dat_data_fp16_16;
reg      [15:0] in_dat_data_fp16_17;
reg      [15:0] in_dat_data_fp16_18;
reg      [15:0] in_dat_data_fp16_19;
reg      [15:0] in_dat_data_fp16_2;
reg      [15:0] in_dat_data_fp16_20;
reg      [15:0] in_dat_data_fp16_21;
reg      [15:0] in_dat_data_fp16_22;
reg      [15:0] in_dat_data_fp16_23;
reg      [15:0] in_dat_data_fp16_24;
reg      [15:0] in_dat_data_fp16_25;
reg      [15:0] in_dat_data_fp16_26;
reg      [15:0] in_dat_data_fp16_27;
reg      [15:0] in_dat_data_fp16_28;
reg      [15:0] in_dat_data_fp16_29;
reg      [15:0] in_dat_data_fp16_3;
reg      [15:0] in_dat_data_fp16_30;
reg      [15:0] in_dat_data_fp16_31;
reg      [15:0] in_dat_data_fp16_32;
reg      [15:0] in_dat_data_fp16_33;
reg      [15:0] in_dat_data_fp16_34;
reg      [15:0] in_dat_data_fp16_35;
reg      [15:0] in_dat_data_fp16_36;
reg      [15:0] in_dat_data_fp16_37;
reg      [15:0] in_dat_data_fp16_38;
reg      [15:0] in_dat_data_fp16_39;
reg      [15:0] in_dat_data_fp16_4;
reg      [15:0] in_dat_data_fp16_40;
reg      [15:0] in_dat_data_fp16_41;
reg      [15:0] in_dat_data_fp16_42;
reg      [15:0] in_dat_data_fp16_43;
reg      [15:0] in_dat_data_fp16_44;
reg      [15:0] in_dat_data_fp16_45;
reg      [15:0] in_dat_data_fp16_46;
reg      [15:0] in_dat_data_fp16_47;
reg      [15:0] in_dat_data_fp16_48;
reg      [15:0] in_dat_data_fp16_49;
reg      [15:0] in_dat_data_fp16_5;
reg      [15:0] in_dat_data_fp16_50;
reg      [15:0] in_dat_data_fp16_51;
reg      [15:0] in_dat_data_fp16_52;
reg      [15:0] in_dat_data_fp16_53;
reg      [15:0] in_dat_data_fp16_54;
reg      [15:0] in_dat_data_fp16_55;
reg      [15:0] in_dat_data_fp16_56;
reg      [15:0] in_dat_data_fp16_57;
reg      [15:0] in_dat_data_fp16_58;
reg      [15:0] in_dat_data_fp16_59;
reg      [15:0] in_dat_data_fp16_6;
reg      [15:0] in_dat_data_fp16_60;
reg      [15:0] in_dat_data_fp16_61;
reg      [15:0] in_dat_data_fp16_62;
reg      [15:0] in_dat_data_fp16_63;
reg      [15:0] in_dat_data_fp16_7;
reg      [15:0] in_dat_data_fp16_8;
reg      [15:0] in_dat_data_fp16_9;
reg      [11:0] in_dat_data_fp16_mts_ori0;
reg      [11:0] in_dat_data_fp16_mts_ori1;
reg      [11:0] in_dat_data_fp16_mts_ori10;
reg      [11:0] in_dat_data_fp16_mts_ori11;
reg      [11:0] in_dat_data_fp16_mts_ori12;
reg      [11:0] in_dat_data_fp16_mts_ori13;
reg      [11:0] in_dat_data_fp16_mts_ori14;
reg      [11:0] in_dat_data_fp16_mts_ori15;
reg      [11:0] in_dat_data_fp16_mts_ori16;
reg      [11:0] in_dat_data_fp16_mts_ori17;
reg      [11:0] in_dat_data_fp16_mts_ori18;
reg      [11:0] in_dat_data_fp16_mts_ori19;
reg      [11:0] in_dat_data_fp16_mts_ori2;
reg      [11:0] in_dat_data_fp16_mts_ori20;
reg      [11:0] in_dat_data_fp16_mts_ori21;
reg      [11:0] in_dat_data_fp16_mts_ori22;
reg      [11:0] in_dat_data_fp16_mts_ori23;
reg      [11:0] in_dat_data_fp16_mts_ori24;
reg      [11:0] in_dat_data_fp16_mts_ori25;
reg      [11:0] in_dat_data_fp16_mts_ori26;
reg      [11:0] in_dat_data_fp16_mts_ori27;
reg      [11:0] in_dat_data_fp16_mts_ori28;
reg      [11:0] in_dat_data_fp16_mts_ori29;
reg      [11:0] in_dat_data_fp16_mts_ori3;
reg      [11:0] in_dat_data_fp16_mts_ori30;
reg      [11:0] in_dat_data_fp16_mts_ori31;
reg      [11:0] in_dat_data_fp16_mts_ori32;
reg      [11:0] in_dat_data_fp16_mts_ori33;
reg      [11:0] in_dat_data_fp16_mts_ori34;
reg      [11:0] in_dat_data_fp16_mts_ori35;
reg      [11:0] in_dat_data_fp16_mts_ori36;
reg      [11:0] in_dat_data_fp16_mts_ori37;
reg      [11:0] in_dat_data_fp16_mts_ori38;
reg      [11:0] in_dat_data_fp16_mts_ori39;
reg      [11:0] in_dat_data_fp16_mts_ori4;
reg      [11:0] in_dat_data_fp16_mts_ori40;
reg      [11:0] in_dat_data_fp16_mts_ori41;
reg      [11:0] in_dat_data_fp16_mts_ori42;
reg      [11:0] in_dat_data_fp16_mts_ori43;
reg      [11:0] in_dat_data_fp16_mts_ori44;
reg      [11:0] in_dat_data_fp16_mts_ori45;
reg      [11:0] in_dat_data_fp16_mts_ori46;
reg      [11:0] in_dat_data_fp16_mts_ori47;
reg      [11:0] in_dat_data_fp16_mts_ori48;
reg      [11:0] in_dat_data_fp16_mts_ori49;
reg      [11:0] in_dat_data_fp16_mts_ori5;
reg      [11:0] in_dat_data_fp16_mts_ori50;
reg      [11:0] in_dat_data_fp16_mts_ori51;
reg      [11:0] in_dat_data_fp16_mts_ori52;
reg      [11:0] in_dat_data_fp16_mts_ori53;
reg      [11:0] in_dat_data_fp16_mts_ori54;
reg      [11:0] in_dat_data_fp16_mts_ori55;
reg      [11:0] in_dat_data_fp16_mts_ori56;
reg      [11:0] in_dat_data_fp16_mts_ori57;
reg      [11:0] in_dat_data_fp16_mts_ori58;
reg      [11:0] in_dat_data_fp16_mts_ori59;
reg      [11:0] in_dat_data_fp16_mts_ori6;
reg      [11:0] in_dat_data_fp16_mts_ori60;
reg      [11:0] in_dat_data_fp16_mts_ori61;
reg      [11:0] in_dat_data_fp16_mts_ori62;
reg      [11:0] in_dat_data_fp16_mts_ori63;
reg      [11:0] in_dat_data_fp16_mts_ori7;
reg      [11:0] in_dat_data_fp16_mts_ori8;
reg      [11:0] in_dat_data_fp16_mts_ori9;
reg      [14:0] in_dat_data_fp16_mts_sft0;
reg      [14:0] in_dat_data_fp16_mts_sft1;
reg      [14:0] in_dat_data_fp16_mts_sft10;
reg      [14:0] in_dat_data_fp16_mts_sft11;
reg      [14:0] in_dat_data_fp16_mts_sft12;
reg      [14:0] in_dat_data_fp16_mts_sft13;
reg      [14:0] in_dat_data_fp16_mts_sft14;
reg      [14:0] in_dat_data_fp16_mts_sft15;
reg      [14:0] in_dat_data_fp16_mts_sft16;
reg      [14:0] in_dat_data_fp16_mts_sft17;
reg      [14:0] in_dat_data_fp16_mts_sft18;
reg      [14:0] in_dat_data_fp16_mts_sft19;
reg      [14:0] in_dat_data_fp16_mts_sft2;
reg      [14:0] in_dat_data_fp16_mts_sft20;
reg      [14:0] in_dat_data_fp16_mts_sft21;
reg      [14:0] in_dat_data_fp16_mts_sft22;
reg      [14:0] in_dat_data_fp16_mts_sft23;
reg      [14:0] in_dat_data_fp16_mts_sft24;
reg      [14:0] in_dat_data_fp16_mts_sft25;
reg      [14:0] in_dat_data_fp16_mts_sft26;
reg      [14:0] in_dat_data_fp16_mts_sft27;
reg      [14:0] in_dat_data_fp16_mts_sft28;
reg      [14:0] in_dat_data_fp16_mts_sft29;
reg      [14:0] in_dat_data_fp16_mts_sft3;
reg      [14:0] in_dat_data_fp16_mts_sft30;
reg      [14:0] in_dat_data_fp16_mts_sft31;
reg      [14:0] in_dat_data_fp16_mts_sft32;
reg      [14:0] in_dat_data_fp16_mts_sft33;
reg      [14:0] in_dat_data_fp16_mts_sft34;
reg      [14:0] in_dat_data_fp16_mts_sft35;
reg      [14:0] in_dat_data_fp16_mts_sft36;
reg      [14:0] in_dat_data_fp16_mts_sft37;
reg      [14:0] in_dat_data_fp16_mts_sft38;
reg      [14:0] in_dat_data_fp16_mts_sft39;
reg      [14:0] in_dat_data_fp16_mts_sft4;
reg      [14:0] in_dat_data_fp16_mts_sft40;
reg      [14:0] in_dat_data_fp16_mts_sft41;
reg      [14:0] in_dat_data_fp16_mts_sft42;
reg      [14:0] in_dat_data_fp16_mts_sft43;
reg      [14:0] in_dat_data_fp16_mts_sft44;
reg      [14:0] in_dat_data_fp16_mts_sft45;
reg      [14:0] in_dat_data_fp16_mts_sft46;
reg      [14:0] in_dat_data_fp16_mts_sft47;
reg      [14:0] in_dat_data_fp16_mts_sft48;
reg      [14:0] in_dat_data_fp16_mts_sft49;
reg      [14:0] in_dat_data_fp16_mts_sft5;
reg      [14:0] in_dat_data_fp16_mts_sft50;
reg      [14:0] in_dat_data_fp16_mts_sft51;
reg      [14:0] in_dat_data_fp16_mts_sft52;
reg      [14:0] in_dat_data_fp16_mts_sft53;
reg      [14:0] in_dat_data_fp16_mts_sft54;
reg      [14:0] in_dat_data_fp16_mts_sft55;
reg      [14:0] in_dat_data_fp16_mts_sft56;
reg      [14:0] in_dat_data_fp16_mts_sft57;
reg      [14:0] in_dat_data_fp16_mts_sft58;
reg      [14:0] in_dat_data_fp16_mts_sft59;
reg      [14:0] in_dat_data_fp16_mts_sft6;
reg      [14:0] in_dat_data_fp16_mts_sft60;
reg      [14:0] in_dat_data_fp16_mts_sft61;
reg      [14:0] in_dat_data_fp16_mts_sft62;
reg      [14:0] in_dat_data_fp16_mts_sft63;
reg      [14:0] in_dat_data_fp16_mts_sft7;
reg      [14:0] in_dat_data_fp16_mts_sft8;
reg      [14:0] in_dat_data_fp16_mts_sft9;
reg    [1023:0] in_dat_data_int16;
reg      [15:0] in_dat_data_int16_0;
reg      [15:0] in_dat_data_int16_1;
reg      [15:0] in_dat_data_int16_10;
reg      [15:0] in_dat_data_int16_11;
reg      [15:0] in_dat_data_int16_12;
reg      [15:0] in_dat_data_int16_13;
reg      [15:0] in_dat_data_int16_14;
reg      [15:0] in_dat_data_int16_15;
reg      [15:0] in_dat_data_int16_16;
reg      [15:0] in_dat_data_int16_17;
reg      [15:0] in_dat_data_int16_18;
reg      [15:0] in_dat_data_int16_19;
reg      [15:0] in_dat_data_int16_2;
reg      [15:0] in_dat_data_int16_20;
reg      [15:0] in_dat_data_int16_21;
reg      [15:0] in_dat_data_int16_22;
reg      [15:0] in_dat_data_int16_23;
reg      [15:0] in_dat_data_int16_24;
reg      [15:0] in_dat_data_int16_25;
reg      [15:0] in_dat_data_int16_26;
reg      [15:0] in_dat_data_int16_27;
reg      [15:0] in_dat_data_int16_28;
reg      [15:0] in_dat_data_int16_29;
reg      [15:0] in_dat_data_int16_3;
reg      [15:0] in_dat_data_int16_30;
reg      [15:0] in_dat_data_int16_31;
reg      [15:0] in_dat_data_int16_32;
reg      [15:0] in_dat_data_int16_33;
reg      [15:0] in_dat_data_int16_34;
reg      [15:0] in_dat_data_int16_35;
reg      [15:0] in_dat_data_int16_36;
reg      [15:0] in_dat_data_int16_37;
reg      [15:0] in_dat_data_int16_38;
reg      [15:0] in_dat_data_int16_39;
reg      [15:0] in_dat_data_int16_4;
reg      [15:0] in_dat_data_int16_40;
reg      [15:0] in_dat_data_int16_41;
reg      [15:0] in_dat_data_int16_42;
reg      [15:0] in_dat_data_int16_43;
reg      [15:0] in_dat_data_int16_44;
reg      [15:0] in_dat_data_int16_45;
reg      [15:0] in_dat_data_int16_46;
reg      [15:0] in_dat_data_int16_47;
reg      [15:0] in_dat_data_int16_48;
reg      [15:0] in_dat_data_int16_49;
reg      [15:0] in_dat_data_int16_5;
reg      [15:0] in_dat_data_int16_50;
reg      [15:0] in_dat_data_int16_51;
reg      [15:0] in_dat_data_int16_52;
reg      [15:0] in_dat_data_int16_53;
reg      [15:0] in_dat_data_int16_54;
reg      [15:0] in_dat_data_int16_55;
reg      [15:0] in_dat_data_int16_56;
reg      [15:0] in_dat_data_int16_57;
reg      [15:0] in_dat_data_int16_58;
reg      [15:0] in_dat_data_int16_59;
reg      [15:0] in_dat_data_int16_6;
reg      [15:0] in_dat_data_int16_60;
reg      [15:0] in_dat_data_int16_61;
reg      [15:0] in_dat_data_int16_62;
reg      [15:0] in_dat_data_int16_63;
reg      [15:0] in_dat_data_int16_7;
reg      [15:0] in_dat_data_int16_8;
reg      [15:0] in_dat_data_int16_9;
reg    [1023:0] in_dat_data_int8;
reg      [15:0] in_dat_data_int8_0;
reg      [15:0] in_dat_data_int8_1;
reg      [15:0] in_dat_data_int8_10;
reg      [15:0] in_dat_data_int8_11;
reg      [15:0] in_dat_data_int8_12;
reg      [15:0] in_dat_data_int8_13;
reg      [15:0] in_dat_data_int8_14;
reg      [15:0] in_dat_data_int8_15;
reg      [15:0] in_dat_data_int8_16;
reg      [15:0] in_dat_data_int8_17;
reg      [15:0] in_dat_data_int8_18;
reg      [15:0] in_dat_data_int8_19;
reg      [15:0] in_dat_data_int8_2;
reg      [15:0] in_dat_data_int8_20;
reg      [15:0] in_dat_data_int8_21;
reg      [15:0] in_dat_data_int8_22;
reg      [15:0] in_dat_data_int8_23;
reg      [15:0] in_dat_data_int8_24;
reg      [15:0] in_dat_data_int8_25;
reg      [15:0] in_dat_data_int8_26;
reg      [15:0] in_dat_data_int8_27;
reg      [15:0] in_dat_data_int8_28;
reg      [15:0] in_dat_data_int8_29;
reg      [15:0] in_dat_data_int8_3;
reg      [15:0] in_dat_data_int8_30;
reg      [15:0] in_dat_data_int8_31;
reg      [15:0] in_dat_data_int8_32;
reg      [15:0] in_dat_data_int8_33;
reg      [15:0] in_dat_data_int8_34;
reg      [15:0] in_dat_data_int8_35;
reg      [15:0] in_dat_data_int8_36;
reg      [15:0] in_dat_data_int8_37;
reg      [15:0] in_dat_data_int8_38;
reg      [15:0] in_dat_data_int8_39;
reg      [15:0] in_dat_data_int8_4;
reg      [15:0] in_dat_data_int8_40;
reg      [15:0] in_dat_data_int8_41;
reg      [15:0] in_dat_data_int8_42;
reg      [15:0] in_dat_data_int8_43;
reg      [15:0] in_dat_data_int8_44;
reg      [15:0] in_dat_data_int8_45;
reg      [15:0] in_dat_data_int8_46;
reg      [15:0] in_dat_data_int8_47;
reg      [15:0] in_dat_data_int8_48;
reg      [15:0] in_dat_data_int8_49;
reg      [15:0] in_dat_data_int8_5;
reg      [15:0] in_dat_data_int8_50;
reg      [15:0] in_dat_data_int8_51;
reg      [15:0] in_dat_data_int8_52;
reg      [15:0] in_dat_data_int8_53;
reg      [15:0] in_dat_data_int8_54;
reg      [15:0] in_dat_data_int8_55;
reg      [15:0] in_dat_data_int8_56;
reg      [15:0] in_dat_data_int8_57;
reg      [15:0] in_dat_data_int8_58;
reg      [15:0] in_dat_data_int8_59;
reg      [15:0] in_dat_data_int8_6;
reg      [15:0] in_dat_data_int8_60;
reg      [15:0] in_dat_data_int8_61;
reg      [15:0] in_dat_data_int8_62;
reg      [15:0] in_dat_data_int8_63;
reg      [15:0] in_dat_data_int8_7;
reg      [15:0] in_dat_data_int8_8;
reg      [15:0] in_dat_data_int8_9;
reg    [1023:0] in_dat_data_pack;
reg     [191:0] in_dat_exp;
reg     [127:0] in_dat_mask_int8;
reg      [63:0] in_dat_nan;
reg      [63:0] in_dat_norm;
reg    [1023:0] in_wt_data_fp16;
reg      [15:0] in_wt_data_fp16_0;
reg      [15:0] in_wt_data_fp16_1;
reg      [15:0] in_wt_data_fp16_10;
reg      [15:0] in_wt_data_fp16_11;
reg      [15:0] in_wt_data_fp16_12;
reg      [15:0] in_wt_data_fp16_13;
reg      [15:0] in_wt_data_fp16_14;
reg      [15:0] in_wt_data_fp16_15;
reg      [15:0] in_wt_data_fp16_16;
reg      [15:0] in_wt_data_fp16_17;
reg      [15:0] in_wt_data_fp16_18;
reg      [15:0] in_wt_data_fp16_19;
reg      [15:0] in_wt_data_fp16_2;
reg      [15:0] in_wt_data_fp16_20;
reg      [15:0] in_wt_data_fp16_21;
reg      [15:0] in_wt_data_fp16_22;
reg      [15:0] in_wt_data_fp16_23;
reg      [15:0] in_wt_data_fp16_24;
reg      [15:0] in_wt_data_fp16_25;
reg      [15:0] in_wt_data_fp16_26;
reg      [15:0] in_wt_data_fp16_27;
reg      [15:0] in_wt_data_fp16_28;
reg      [15:0] in_wt_data_fp16_29;
reg      [15:0] in_wt_data_fp16_3;
reg      [15:0] in_wt_data_fp16_30;
reg      [15:0] in_wt_data_fp16_31;
reg      [15:0] in_wt_data_fp16_32;
reg      [15:0] in_wt_data_fp16_33;
reg      [15:0] in_wt_data_fp16_34;
reg      [15:0] in_wt_data_fp16_35;
reg      [15:0] in_wt_data_fp16_36;
reg      [15:0] in_wt_data_fp16_37;
reg      [15:0] in_wt_data_fp16_38;
reg      [15:0] in_wt_data_fp16_39;
reg      [15:0] in_wt_data_fp16_4;
reg      [15:0] in_wt_data_fp16_40;
reg      [15:0] in_wt_data_fp16_41;
reg      [15:0] in_wt_data_fp16_42;
reg      [15:0] in_wt_data_fp16_43;
reg      [15:0] in_wt_data_fp16_44;
reg      [15:0] in_wt_data_fp16_45;
reg      [15:0] in_wt_data_fp16_46;
reg      [15:0] in_wt_data_fp16_47;
reg      [15:0] in_wt_data_fp16_48;
reg      [15:0] in_wt_data_fp16_49;
reg      [15:0] in_wt_data_fp16_5;
reg      [15:0] in_wt_data_fp16_50;
reg      [15:0] in_wt_data_fp16_51;
reg      [15:0] in_wt_data_fp16_52;
reg      [15:0] in_wt_data_fp16_53;
reg      [15:0] in_wt_data_fp16_54;
reg      [15:0] in_wt_data_fp16_55;
reg      [15:0] in_wt_data_fp16_56;
reg      [15:0] in_wt_data_fp16_57;
reg      [15:0] in_wt_data_fp16_58;
reg      [15:0] in_wt_data_fp16_59;
reg      [15:0] in_wt_data_fp16_6;
reg      [15:0] in_wt_data_fp16_60;
reg      [15:0] in_wt_data_fp16_61;
reg      [15:0] in_wt_data_fp16_62;
reg      [15:0] in_wt_data_fp16_63;
reg      [15:0] in_wt_data_fp16_7;
reg      [15:0] in_wt_data_fp16_8;
reg      [15:0] in_wt_data_fp16_9;
reg      [11:0] in_wt_data_fp16_mts_ori0;
reg      [11:0] in_wt_data_fp16_mts_ori1;
reg      [11:0] in_wt_data_fp16_mts_ori10;
reg      [11:0] in_wt_data_fp16_mts_ori11;
reg      [11:0] in_wt_data_fp16_mts_ori12;
reg      [11:0] in_wt_data_fp16_mts_ori13;
reg      [11:0] in_wt_data_fp16_mts_ori14;
reg      [11:0] in_wt_data_fp16_mts_ori15;
reg      [11:0] in_wt_data_fp16_mts_ori16;
reg      [11:0] in_wt_data_fp16_mts_ori17;
reg      [11:0] in_wt_data_fp16_mts_ori18;
reg      [11:0] in_wt_data_fp16_mts_ori19;
reg      [11:0] in_wt_data_fp16_mts_ori2;
reg      [11:0] in_wt_data_fp16_mts_ori20;
reg      [11:0] in_wt_data_fp16_mts_ori21;
reg      [11:0] in_wt_data_fp16_mts_ori22;
reg      [11:0] in_wt_data_fp16_mts_ori23;
reg      [11:0] in_wt_data_fp16_mts_ori24;
reg      [11:0] in_wt_data_fp16_mts_ori25;
reg      [11:0] in_wt_data_fp16_mts_ori26;
reg      [11:0] in_wt_data_fp16_mts_ori27;
reg      [11:0] in_wt_data_fp16_mts_ori28;
reg      [11:0] in_wt_data_fp16_mts_ori29;
reg      [11:0] in_wt_data_fp16_mts_ori3;
reg      [11:0] in_wt_data_fp16_mts_ori30;
reg      [11:0] in_wt_data_fp16_mts_ori31;
reg      [11:0] in_wt_data_fp16_mts_ori32;
reg      [11:0] in_wt_data_fp16_mts_ori33;
reg      [11:0] in_wt_data_fp16_mts_ori34;
reg      [11:0] in_wt_data_fp16_mts_ori35;
reg      [11:0] in_wt_data_fp16_mts_ori36;
reg      [11:0] in_wt_data_fp16_mts_ori37;
reg      [11:0] in_wt_data_fp16_mts_ori38;
reg      [11:0] in_wt_data_fp16_mts_ori39;
reg      [11:0] in_wt_data_fp16_mts_ori4;
reg      [11:0] in_wt_data_fp16_mts_ori40;
reg      [11:0] in_wt_data_fp16_mts_ori41;
reg      [11:0] in_wt_data_fp16_mts_ori42;
reg      [11:0] in_wt_data_fp16_mts_ori43;
reg      [11:0] in_wt_data_fp16_mts_ori44;
reg      [11:0] in_wt_data_fp16_mts_ori45;
reg      [11:0] in_wt_data_fp16_mts_ori46;
reg      [11:0] in_wt_data_fp16_mts_ori47;
reg      [11:0] in_wt_data_fp16_mts_ori48;
reg      [11:0] in_wt_data_fp16_mts_ori49;
reg      [11:0] in_wt_data_fp16_mts_ori5;
reg      [11:0] in_wt_data_fp16_mts_ori50;
reg      [11:0] in_wt_data_fp16_mts_ori51;
reg      [11:0] in_wt_data_fp16_mts_ori52;
reg      [11:0] in_wt_data_fp16_mts_ori53;
reg      [11:0] in_wt_data_fp16_mts_ori54;
reg      [11:0] in_wt_data_fp16_mts_ori55;
reg      [11:0] in_wt_data_fp16_mts_ori56;
reg      [11:0] in_wt_data_fp16_mts_ori57;
reg      [11:0] in_wt_data_fp16_mts_ori58;
reg      [11:0] in_wt_data_fp16_mts_ori59;
reg      [11:0] in_wt_data_fp16_mts_ori6;
reg      [11:0] in_wt_data_fp16_mts_ori60;
reg      [11:0] in_wt_data_fp16_mts_ori61;
reg      [11:0] in_wt_data_fp16_mts_ori62;
reg      [11:0] in_wt_data_fp16_mts_ori63;
reg      [11:0] in_wt_data_fp16_mts_ori7;
reg      [11:0] in_wt_data_fp16_mts_ori8;
reg      [11:0] in_wt_data_fp16_mts_ori9;
reg      [14:0] in_wt_data_fp16_mts_sft0;
reg      [14:0] in_wt_data_fp16_mts_sft1;
reg      [14:0] in_wt_data_fp16_mts_sft10;
reg      [14:0] in_wt_data_fp16_mts_sft11;
reg      [14:0] in_wt_data_fp16_mts_sft12;
reg      [14:0] in_wt_data_fp16_mts_sft13;
reg      [14:0] in_wt_data_fp16_mts_sft14;
reg      [14:0] in_wt_data_fp16_mts_sft15;
reg      [14:0] in_wt_data_fp16_mts_sft16;
reg      [14:0] in_wt_data_fp16_mts_sft17;
reg      [14:0] in_wt_data_fp16_mts_sft18;
reg      [14:0] in_wt_data_fp16_mts_sft19;
reg      [14:0] in_wt_data_fp16_mts_sft2;
reg      [14:0] in_wt_data_fp16_mts_sft20;
reg      [14:0] in_wt_data_fp16_mts_sft21;
reg      [14:0] in_wt_data_fp16_mts_sft22;
reg      [14:0] in_wt_data_fp16_mts_sft23;
reg      [14:0] in_wt_data_fp16_mts_sft24;
reg      [14:0] in_wt_data_fp16_mts_sft25;
reg      [14:0] in_wt_data_fp16_mts_sft26;
reg      [14:0] in_wt_data_fp16_mts_sft27;
reg      [14:0] in_wt_data_fp16_mts_sft28;
reg      [14:0] in_wt_data_fp16_mts_sft29;
reg      [14:0] in_wt_data_fp16_mts_sft3;
reg      [14:0] in_wt_data_fp16_mts_sft30;
reg      [14:0] in_wt_data_fp16_mts_sft31;
reg      [14:0] in_wt_data_fp16_mts_sft32;
reg      [14:0] in_wt_data_fp16_mts_sft33;
reg      [14:0] in_wt_data_fp16_mts_sft34;
reg      [14:0] in_wt_data_fp16_mts_sft35;
reg      [14:0] in_wt_data_fp16_mts_sft36;
reg      [14:0] in_wt_data_fp16_mts_sft37;
reg      [14:0] in_wt_data_fp16_mts_sft38;
reg      [14:0] in_wt_data_fp16_mts_sft39;
reg      [14:0] in_wt_data_fp16_mts_sft4;
reg      [14:0] in_wt_data_fp16_mts_sft40;
reg      [14:0] in_wt_data_fp16_mts_sft41;
reg      [14:0] in_wt_data_fp16_mts_sft42;
reg      [14:0] in_wt_data_fp16_mts_sft43;
reg      [14:0] in_wt_data_fp16_mts_sft44;
reg      [14:0] in_wt_data_fp16_mts_sft45;
reg      [14:0] in_wt_data_fp16_mts_sft46;
reg      [14:0] in_wt_data_fp16_mts_sft47;
reg      [14:0] in_wt_data_fp16_mts_sft48;
reg      [14:0] in_wt_data_fp16_mts_sft49;
reg      [14:0] in_wt_data_fp16_mts_sft5;
reg      [14:0] in_wt_data_fp16_mts_sft50;
reg      [14:0] in_wt_data_fp16_mts_sft51;
reg      [14:0] in_wt_data_fp16_mts_sft52;
reg      [14:0] in_wt_data_fp16_mts_sft53;
reg      [14:0] in_wt_data_fp16_mts_sft54;
reg      [14:0] in_wt_data_fp16_mts_sft55;
reg      [14:0] in_wt_data_fp16_mts_sft56;
reg      [14:0] in_wt_data_fp16_mts_sft57;
reg      [14:0] in_wt_data_fp16_mts_sft58;
reg      [14:0] in_wt_data_fp16_mts_sft59;
reg      [14:0] in_wt_data_fp16_mts_sft6;
reg      [14:0] in_wt_data_fp16_mts_sft60;
reg      [14:0] in_wt_data_fp16_mts_sft61;
reg      [14:0] in_wt_data_fp16_mts_sft62;
reg      [14:0] in_wt_data_fp16_mts_sft63;
reg      [14:0] in_wt_data_fp16_mts_sft7;
reg      [14:0] in_wt_data_fp16_mts_sft8;
reg      [14:0] in_wt_data_fp16_mts_sft9;
reg    [1023:0] in_wt_data_int16;
reg      [15:0] in_wt_data_int16_0;
reg      [15:0] in_wt_data_int16_1;
reg      [15:0] in_wt_data_int16_10;
reg      [15:0] in_wt_data_int16_11;
reg      [15:0] in_wt_data_int16_12;
reg      [15:0] in_wt_data_int16_13;
reg      [15:0] in_wt_data_int16_14;
reg      [15:0] in_wt_data_int16_15;
reg      [15:0] in_wt_data_int16_16;
reg      [15:0] in_wt_data_int16_17;
reg      [15:0] in_wt_data_int16_18;
reg      [15:0] in_wt_data_int16_19;
reg      [15:0] in_wt_data_int16_2;
reg      [15:0] in_wt_data_int16_20;
reg      [15:0] in_wt_data_int16_21;
reg      [15:0] in_wt_data_int16_22;
reg      [15:0] in_wt_data_int16_23;
reg      [15:0] in_wt_data_int16_24;
reg      [15:0] in_wt_data_int16_25;
reg      [15:0] in_wt_data_int16_26;
reg      [15:0] in_wt_data_int16_27;
reg      [15:0] in_wt_data_int16_28;
reg      [15:0] in_wt_data_int16_29;
reg      [15:0] in_wt_data_int16_3;
reg      [15:0] in_wt_data_int16_30;
reg      [15:0] in_wt_data_int16_31;
reg      [15:0] in_wt_data_int16_32;
reg      [15:0] in_wt_data_int16_33;
reg      [15:0] in_wt_data_int16_34;
reg      [15:0] in_wt_data_int16_35;
reg      [15:0] in_wt_data_int16_36;
reg      [15:0] in_wt_data_int16_37;
reg      [15:0] in_wt_data_int16_38;
reg      [15:0] in_wt_data_int16_39;
reg      [15:0] in_wt_data_int16_4;
reg      [15:0] in_wt_data_int16_40;
reg      [15:0] in_wt_data_int16_41;
reg      [15:0] in_wt_data_int16_42;
reg      [15:0] in_wt_data_int16_43;
reg      [15:0] in_wt_data_int16_44;
reg      [15:0] in_wt_data_int16_45;
reg      [15:0] in_wt_data_int16_46;
reg      [15:0] in_wt_data_int16_47;
reg      [15:0] in_wt_data_int16_48;
reg      [15:0] in_wt_data_int16_49;
reg      [15:0] in_wt_data_int16_5;
reg      [15:0] in_wt_data_int16_50;
reg      [15:0] in_wt_data_int16_51;
reg      [15:0] in_wt_data_int16_52;
reg      [15:0] in_wt_data_int16_53;
reg      [15:0] in_wt_data_int16_54;
reg      [15:0] in_wt_data_int16_55;
reg      [15:0] in_wt_data_int16_56;
reg      [15:0] in_wt_data_int16_57;
reg      [15:0] in_wt_data_int16_58;
reg      [15:0] in_wt_data_int16_59;
reg      [15:0] in_wt_data_int16_6;
reg      [15:0] in_wt_data_int16_60;
reg      [15:0] in_wt_data_int16_61;
reg      [15:0] in_wt_data_int16_62;
reg      [15:0] in_wt_data_int16_63;
reg      [15:0] in_wt_data_int16_7;
reg      [15:0] in_wt_data_int16_8;
reg      [15:0] in_wt_data_int16_9;
reg    [1023:0] in_wt_data_int8;
reg      [15:0] in_wt_data_int8_0;
reg      [15:0] in_wt_data_int8_1;
reg      [15:0] in_wt_data_int8_10;
reg      [15:0] in_wt_data_int8_11;
reg      [15:0] in_wt_data_int8_12;
reg      [15:0] in_wt_data_int8_13;
reg      [15:0] in_wt_data_int8_14;
reg      [15:0] in_wt_data_int8_15;
reg      [15:0] in_wt_data_int8_16;
reg      [15:0] in_wt_data_int8_17;
reg      [15:0] in_wt_data_int8_18;
reg      [15:0] in_wt_data_int8_19;
reg      [15:0] in_wt_data_int8_2;
reg      [15:0] in_wt_data_int8_20;
reg      [15:0] in_wt_data_int8_21;
reg      [15:0] in_wt_data_int8_22;
reg      [15:0] in_wt_data_int8_23;
reg      [15:0] in_wt_data_int8_24;
reg      [15:0] in_wt_data_int8_25;
reg      [15:0] in_wt_data_int8_26;
reg      [15:0] in_wt_data_int8_27;
reg      [15:0] in_wt_data_int8_28;
reg      [15:0] in_wt_data_int8_29;
reg      [15:0] in_wt_data_int8_3;
reg      [15:0] in_wt_data_int8_30;
reg      [15:0] in_wt_data_int8_31;
reg      [15:0] in_wt_data_int8_32;
reg      [15:0] in_wt_data_int8_33;
reg      [15:0] in_wt_data_int8_34;
reg      [15:0] in_wt_data_int8_35;
reg      [15:0] in_wt_data_int8_36;
reg      [15:0] in_wt_data_int8_37;
reg      [15:0] in_wt_data_int8_38;
reg      [15:0] in_wt_data_int8_39;
reg      [15:0] in_wt_data_int8_4;
reg      [15:0] in_wt_data_int8_40;
reg      [15:0] in_wt_data_int8_41;
reg      [15:0] in_wt_data_int8_42;
reg      [15:0] in_wt_data_int8_43;
reg      [15:0] in_wt_data_int8_44;
reg      [15:0] in_wt_data_int8_45;
reg      [15:0] in_wt_data_int8_46;
reg      [15:0] in_wt_data_int8_47;
reg      [15:0] in_wt_data_int8_48;
reg      [15:0] in_wt_data_int8_49;
reg      [15:0] in_wt_data_int8_5;
reg      [15:0] in_wt_data_int8_50;
reg      [15:0] in_wt_data_int8_51;
reg      [15:0] in_wt_data_int8_52;
reg      [15:0] in_wt_data_int8_53;
reg      [15:0] in_wt_data_int8_54;
reg      [15:0] in_wt_data_int8_55;
reg      [15:0] in_wt_data_int8_56;
reg      [15:0] in_wt_data_int8_57;
reg      [15:0] in_wt_data_int8_58;
reg      [15:0] in_wt_data_int8_59;
reg      [15:0] in_wt_data_int8_6;
reg      [15:0] in_wt_data_int8_60;
reg      [15:0] in_wt_data_int8_61;
reg      [15:0] in_wt_data_int8_62;
reg      [15:0] in_wt_data_int8_63;
reg      [15:0] in_wt_data_int8_7;
reg      [15:0] in_wt_data_int8_8;
reg      [15:0] in_wt_data_int8_9;
reg    [1023:0] in_wt_data_pack;
reg     [191:0] in_wt_exp;
reg     [127:0] in_wt_mask_int8;
reg      [63:0] in_wt_nan;
reg      [63:0] in_wt_norm;
reg    [1023:0] wt0_actv_data;
reg      [63:0] wt0_actv_nan;
reg     [127:0] wt0_actv_nz;
reg     [103:0] wt0_actv_pvld;
reg             wt0_actv_pvld_w;
reg       [0:0] wt0_actv_vld;
reg    [1023:0] wt0_sd_data;
reg     [191:0] wt0_sd_exp;
reg      [63:0] wt0_sd_mask;
reg      [63:0] wt0_sd_nan;
reg     [127:0] wt0_sd_nz;
reg             wt0_sd_pvld;
reg             wt0_sd_pvld_w;
reg    [1023:0] wt1_actv_data;
reg      [63:0] wt1_actv_nan;
reg     [127:0] wt1_actv_nz;
reg     [103:0] wt1_actv_pvld;
reg             wt1_actv_pvld_w;
reg       [0:0] wt1_actv_vld;
reg    [1023:0] wt1_sd_data;
reg     [191:0] wt1_sd_exp;
reg      [63:0] wt1_sd_mask;
reg      [63:0] wt1_sd_nan;
reg     [127:0] wt1_sd_nz;
reg             wt1_sd_pvld;
reg             wt1_sd_pvld_w;
reg    [1023:0] wt2_actv_data;
reg      [63:0] wt2_actv_nan;
reg     [127:0] wt2_actv_nz;
reg     [103:0] wt2_actv_pvld;
reg             wt2_actv_pvld_w;
reg       [0:0] wt2_actv_vld;
reg    [1023:0] wt2_sd_data;
reg     [191:0] wt2_sd_exp;
reg      [63:0] wt2_sd_mask;
reg      [63:0] wt2_sd_nan;
reg     [127:0] wt2_sd_nz;
reg             wt2_sd_pvld;
reg             wt2_sd_pvld_w;
reg    [1023:0] wt3_actv_data;
reg      [63:0] wt3_actv_nan;
reg     [127:0] wt3_actv_nz;
reg     [103:0] wt3_actv_pvld;
reg             wt3_actv_pvld_w;
reg       [0:0] wt3_actv_vld;
reg    [1023:0] wt3_sd_data;
reg     [191:0] wt3_sd_exp;
reg      [63:0] wt3_sd_mask;
reg      [63:0] wt3_sd_nan;
reg     [127:0] wt3_sd_nz;
reg             wt3_sd_pvld;
reg             wt3_sd_pvld_w;
reg    [1023:0] wt4_actv_data;
reg      [63:0] wt4_actv_nan;
reg     [127:0] wt4_actv_nz;
reg     [103:0] wt4_actv_pvld;
reg             wt4_actv_pvld_w;
reg       [0:0] wt4_actv_vld;
reg    [1023:0] wt4_sd_data;
reg     [191:0] wt4_sd_exp;
reg      [63:0] wt4_sd_mask;
reg      [63:0] wt4_sd_nan;
reg     [127:0] wt4_sd_nz;
reg             wt4_sd_pvld;
reg             wt4_sd_pvld_w;
reg    [1023:0] wt5_actv_data;
reg      [63:0] wt5_actv_nan;
reg     [127:0] wt5_actv_nz;
reg     [103:0] wt5_actv_pvld;
reg             wt5_actv_pvld_w;
reg       [0:0] wt5_actv_vld;
reg    [1023:0] wt5_sd_data;
reg     [191:0] wt5_sd_exp;
reg      [63:0] wt5_sd_mask;
reg      [63:0] wt5_sd_nan;
reg     [127:0] wt5_sd_nz;
reg             wt5_sd_pvld;
reg             wt5_sd_pvld_w;
reg    [1023:0] wt6_actv_data;
reg      [63:0] wt6_actv_nan;
reg     [127:0] wt6_actv_nz;
reg     [103:0] wt6_actv_pvld;
reg             wt6_actv_pvld_w;
reg       [0:0] wt6_actv_vld;
reg    [1023:0] wt6_sd_data;
reg     [191:0] wt6_sd_exp;
reg      [63:0] wt6_sd_mask;
reg      [63:0] wt6_sd_nan;
reg     [127:0] wt6_sd_nz;
reg             wt6_sd_pvld;
reg             wt6_sd_pvld_w;
reg    [1023:0] wt7_actv_data;
reg      [63:0] wt7_actv_nan;
reg     [127:0] wt7_actv_nz;
reg     [103:0] wt7_actv_pvld;
reg             wt7_actv_pvld_w;
reg       [0:0] wt7_actv_vld;
reg    [1023:0] wt7_sd_data;
reg     [191:0] wt7_sd_exp;
reg      [63:0] wt7_sd_mask;
reg      [63:0] wt7_sd_nan;
reg     [127:0] wt7_sd_nz;
reg             wt7_sd_pvld;
reg             wt7_sd_pvld_w;
reg             wt_has_nan;
reg    [1023:0] wt_pre_data;
reg    [1023:0] wt_pre_data_w;
reg     [191:0] wt_pre_exp;
reg     [191:0] wt_pre_exp_w;
reg      [63:0] wt_pre_mask;
reg      [63:0] wt_pre_mask_w;
reg      [63:0] wt_pre_nan;
reg     [127:0] wt_pre_nz;
reg     [127:0] wt_pre_nz_w;
reg       [7:0] wt_pre_sel;

// synoff nets

// monitor nets

// debug nets

// tie high nets

// tie low nets

// no connect nets

// not all bits used nets

// todo nets

    

//==========================================================
// Input config
//==========================================================

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    cfg_is_int8_d1 <= {65{1'b0}};
  end else begin
  if ((cfg_reg_en) == 1'b1) begin
    cfg_is_int8_d1 <= {65{cfg_is_int8}};
  // VCS coverage off
  end else if ((cfg_reg_en) == 1'b0) begin
  end else begin
    cfg_is_int8_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
  end
end
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_no_x #(0,1,0,"No X's allowed on control signals")      zzz_assert_no_x_1x (nvdla_core_clk, `ASSERT_RESET, 1'd1,  (^(cfg_reg_en))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    cfg_is_fp16_d1 <= {98{1'b0}};
  end else begin
  if ((cfg_reg_en) == 1'b1) begin
    cfg_is_fp16_d1 <= {98{cfg_is_fp16}};
  // VCS coverage off
  end else if ((cfg_reg_en) == 1'b0) begin
  end else begin
    cfg_is_fp16_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
  end
end
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_no_x #(0,1,0,"No X's allowed on control signals")      zzz_assert_no_x_2x (nvdla_core_clk, `ASSERT_RESET, 1'd1,  (^(cfg_reg_en))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    cfg_is_int16_d1 <= {64{1'b0}};
  end else begin
  if ((cfg_reg_en) == 1'b1) begin
    cfg_is_int16_d1 <= {64{cfg_is_int16}};
  // VCS coverage off
  end else if ((cfg_reg_en) == 1'b0) begin
  end else begin
    cfg_is_int16_d1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
  end
end
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_no_x #(0,1,0,"No X's allowed on control signals")      zzz_assert_no_x_3x (nvdla_core_clk, `ASSERT_RESET, 1'd1,  (^(cfg_reg_en))); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON

//==========================================================
// Weight reordering and detect
//==========================================================

always @(
  in_wt_data127
  or in_wt_data126
  or in_wt_data125
  or in_wt_data124
  or in_wt_data123
  or in_wt_data122
  or in_wt_data121
  or in_wt_data120
  or in_wt_data119
  or in_wt_data118
  or in_wt_data117
  or in_wt_data116
  or in_wt_data115
  or in_wt_data114
  or in_wt_data113
  or in_wt_data112
  or in_wt_data111
  or in_wt_data110
  or in_wt_data109
  or in_wt_data108
  or in_wt_data107
  or in_wt_data106
  or in_wt_data105
  or in_wt_data104
  or in_wt_data103
  or in_wt_data102
  or in_wt_data101
  or in_wt_data100
  or in_wt_data99
  or in_wt_data98
  or in_wt_data97
  or in_wt_data96
  or in_wt_data95
  or in_wt_data94
  or in_wt_data93
  or in_wt_data92
  or in_wt_data91
  or in_wt_data90
  or in_wt_data89
  or in_wt_data88
  or in_wt_data87
  or in_wt_data86
  or in_wt_data85
  or in_wt_data84
  or in_wt_data83
  or in_wt_data82
  or in_wt_data81
  or in_wt_data80
  or in_wt_data79
  or in_wt_data78
  or in_wt_data77
  or in_wt_data76
  or in_wt_data75
  or in_wt_data74
  or in_wt_data73
  or in_wt_data72
  or in_wt_data71
  or in_wt_data70
  or in_wt_data69
  or in_wt_data68
  or in_wt_data67
  or in_wt_data66
  or in_wt_data65
  or in_wt_data64
  or in_wt_data63
  or in_wt_data62
  or in_wt_data61
  or in_wt_data60
  or in_wt_data59
  or in_wt_data58
  or in_wt_data57
  or in_wt_data56
  or in_wt_data55
  or in_wt_data54
  or in_wt_data53
  or in_wt_data52
  or in_wt_data51
  or in_wt_data50
  or in_wt_data49
  or in_wt_data48
  or in_wt_data47
  or in_wt_data46
  or in_wt_data45
  or in_wt_data44
  or in_wt_data43
  or in_wt_data42
  or in_wt_data41
  or in_wt_data40
  or in_wt_data39
  or in_wt_data38
  or in_wt_data37
  or in_wt_data36
  or in_wt_data35
  or in_wt_data34
  or in_wt_data33
  or in_wt_data32
  or in_wt_data31
  or in_wt_data30
  or in_wt_data29
  or in_wt_data28
  or in_wt_data27
  or in_wt_data26
  or in_wt_data25
  or in_wt_data24
  or in_wt_data23
  or in_wt_data22
  or in_wt_data21
  or in_wt_data20
  or in_wt_data19
  or in_wt_data18
  or in_wt_data17
  or in_wt_data16
  or in_wt_data15
  or in_wt_data14
  or in_wt_data13
  or in_wt_data12
  or in_wt_data11
  or in_wt_data10
  or in_wt_data9
  or in_wt_data8
  or in_wt_data7
  or in_wt_data6
  or in_wt_data5
  or in_wt_data4
  or in_wt_data3
  or in_wt_data2
  or in_wt_data1
  or in_wt_data0
  ) begin
    in_wt_data_pack = {in_wt_data127, in_wt_data126, in_wt_data125, in_wt_data124, in_wt_data123, in_wt_data122, in_wt_data121, in_wt_data120, in_wt_data119, in_wt_data118, in_wt_data117, in_wt_data116, in_wt_data115, in_wt_data114, in_wt_data113, in_wt_data112, in_wt_data111, in_wt_data110, in_wt_data109, in_wt_data108, in_wt_data107, in_wt_data106, in_wt_data105, in_wt_data104, in_wt_data103, in_wt_data102, in_wt_data101, in_wt_data100, in_wt_data99, in_wt_data98, in_wt_data97, in_wt_data96, in_wt_data95, in_wt_data94, in_wt_data93, in_wt_data92, in_wt_data91, in_wt_data90, in_wt_data89, in_wt_data88, in_wt_data87, in_wt_data86, in_wt_data85, in_wt_data84, in_wt_data83, in_wt_data82, in_wt_data81, in_wt_data80, in_wt_data79, in_wt_data78, in_wt_data77, in_wt_data76, in_wt_data75, in_wt_data74, in_wt_data73, in_wt_data72, in_wt_data71, in_wt_data70, in_wt_data69, in_wt_data68, in_wt_data67, in_wt_data66, in_wt_data65, in_wt_data64, in_wt_data63, in_wt_data62, in_wt_data61, in_wt_data60, in_wt_data59, in_wt_data58, in_wt_data57, in_wt_data56, in_wt_data55, in_wt_data54, in_wt_data53, in_wt_data52, in_wt_data51, in_wt_data50, in_wt_data49, in_wt_data48, in_wt_data47, in_wt_data46, in_wt_data45, in_wt_data44, in_wt_data43, in_wt_data42, in_wt_data41, in_wt_data40, in_wt_data39, in_wt_data38, in_wt_data37, in_wt_data36, in_wt_data35, in_wt_data34, in_wt_data33, in_wt_data32, in_wt_data31, in_wt_data30, in_wt_data29, in_wt_data28, in_wt_data27, in_wt_data26, in_wt_data25, in_wt_data24, in_wt_data23, in_wt_data22, in_wt_data21, in_wt_data20, in_wt_data19, in_wt_data18, in_wt_data17, in_wt_data16, in_wt_data15, in_wt_data14, in_wt_data13, in_wt_data12, in_wt_data11, in_wt_data10, in_wt_data9, in_wt_data8, in_wt_data7, in_wt_data6, in_wt_data5, in_wt_data4, in_wt_data3, in_wt_data2, in_wt_data1, in_wt_data0};
end

//////////////// in_wt_data_int16 ////////////////
always @(
  cfg_is_int16_d1
  or in_wt_data127
  or in_wt_data126
  or in_wt_data125
  or in_wt_data124
  or in_wt_data123
  or in_wt_data122
  or in_wt_data121
  or in_wt_data120
  or in_wt_data119
  or in_wt_data118
  or in_wt_data117
  or in_wt_data116
  or in_wt_data115
  or in_wt_data114
  or in_wt_data113
  or in_wt_data112
  or in_wt_data111
  or in_wt_data110
  or in_wt_data109
  or in_wt_data108
  or in_wt_data107
  or in_wt_data106
  or in_wt_data105
  or in_wt_data104
  or in_wt_data103
  or in_wt_data102
  or in_wt_data101
  or in_wt_data100
  or in_wt_data99
  or in_wt_data98
  or in_wt_data97
  or in_wt_data96
  or in_wt_data95
  or in_wt_data94
  or in_wt_data93
  or in_wt_data92
  or in_wt_data91
  or in_wt_data90
  or in_wt_data89
  or in_wt_data88
  or in_wt_data87
  or in_wt_data86
  or in_wt_data85
  or in_wt_data84
  or in_wt_data83
  or in_wt_data82
  or in_wt_data81
  or in_wt_data80
  or in_wt_data79
  or in_wt_data78
  or in_wt_data77
  or in_wt_data76
  or in_wt_data75
  or in_wt_data74
  or in_wt_data73
  or in_wt_data72
  or in_wt_data71
  or in_wt_data70
  or in_wt_data69
  or in_wt_data68
  or in_wt_data67
  or in_wt_data66
  or in_wt_data65
  or in_wt_data64
  or in_wt_data63
  or in_wt_data62
  or in_wt_data61
  or in_wt_data60
  or in_wt_data59
  or in_wt_data58
  or in_wt_data57
  or in_wt_data56
  or in_wt_data55
  or in_wt_data54
  or in_wt_data53
  or in_wt_data52
  or in_wt_data51
  or in_wt_data50
  or in_wt_data49
  or in_wt_data48
  or in_wt_data47
  or in_wt_data46
  or in_wt_data45
  or in_wt_data44
  or in_wt_data43
  or in_wt_data42
  or in_wt_data41
  or in_wt_data40
  or in_wt_data39
  or in_wt_data38
  or in_wt_data37
  or in_wt_data36
  or in_wt_data35
  or in_wt_data34
  or in_wt_data33
  or in_wt_data32
  or in_wt_data31
  or in_wt_data30
  or in_wt_data29
  or in_wt_data28
  or in_wt_data27
  or in_wt_data26
  or in_wt_data25
  or in_wt_data24
  or in_wt_data23
  or in_wt_data22
  or in_wt_data21
  or in_wt_data20
  or in_wt_data19
  or in_wt_data18
  or in_wt_data17
  or in_wt_data16
  or in_wt_data15
  or in_wt_data14
  or in_wt_data13
  or in_wt_data12
  or in_wt_data11
  or in_wt_data10
  or in_wt_data9
  or in_wt_data8
  or in_wt_data7
  or in_wt_data6
  or in_wt_data5
  or in_wt_data4
  or in_wt_data3
  or in_wt_data2
  or in_wt_data1
  or in_wt_data0
  ) begin
    in_wt_data_int16_63 = ({16{cfg_is_int16_d1[63]}} & {in_wt_data127, in_wt_data126});
    in_wt_data_int16_62 = ({16{cfg_is_int16_d1[62]}} & {in_wt_data125, in_wt_data124});
    in_wt_data_int16_61 = ({16{cfg_is_int16_d1[61]}} & {in_wt_data123, in_wt_data122});
    in_wt_data_int16_60 = ({16{cfg_is_int16_d1[60]}} & {in_wt_data121, in_wt_data120});
    in_wt_data_int16_59 = ({16{cfg_is_int16_d1[59]}} & {in_wt_data119, in_wt_data118});
    in_wt_data_int16_58 = ({16{cfg_is_int16_d1[58]}} & {in_wt_data117, in_wt_data116});
    in_wt_data_int16_57 = ({16{cfg_is_int16_d1[57]}} & {in_wt_data115, in_wt_data114});
    in_wt_data_int16_56 = ({16{cfg_is_int16_d1[56]}} & {in_wt_data113, in_wt_data112});
    in_wt_data_int16_55 = ({16{cfg_is_int16_d1[55]}} & {in_wt_data111, in_wt_data110});
    in_wt_data_int16_54 = ({16{cfg_is_int16_d1[54]}} & {in_wt_data109, in_wt_data108});
    in_wt_data_int16_53 = ({16{cfg_is_int16_d1[53]}} & {in_wt_data107, in_wt_data106});
    in_wt_data_int16_52 = ({16{cfg_is_int16_d1[52]}} & {in_wt_data105, in_wt_data104});
    in_wt_data_int16_51 = ({16{cfg_is_int16_d1[51]}} & {in_wt_data103, in_wt_data102});
    in_wt_data_int16_50 = ({16{cfg_is_int16_d1[50]}} & {in_wt_data101, in_wt_data100});
    in_wt_data_int16_49 = ({16{cfg_is_int16_d1[49]}} & {in_wt_data99, in_wt_data98});
    in_wt_data_int16_48 = ({16{cfg_is_int16_d1[48]}} & {in_wt_data97, in_wt_data96});
    in_wt_data_int16_47 = ({16{cfg_is_int16_d1[47]}} & {in_wt_data95, in_wt_data94});
    in_wt_data_int16_46 = ({16{cfg_is_int16_d1[46]}} & {in_wt_data93, in_wt_data92});
    in_wt_data_int16_45 = ({16{cfg_is_int16_d1[45]}} & {in_wt_data91, in_wt_data90});
    in_wt_data_int16_44 = ({16{cfg_is_int16_d1[44]}} & {in_wt_data89, in_wt_data88});
    in_wt_data_int16_43 = ({16{cfg_is_int16_d1[43]}} & {in_wt_data87, in_wt_data86});
    in_wt_data_int16_42 = ({16{cfg_is_int16_d1[42]}} & {in_wt_data85, in_wt_data84});
    in_wt_data_int16_41 = ({16{cfg_is_int16_d1[41]}} & {in_wt_data83, in_wt_data82});
    in_wt_data_int16_40 = ({16{cfg_is_int16_d1[40]}} & {in_wt_data81, in_wt_data80});
    in_wt_data_int16_39 = ({16{cfg_is_int16_d1[39]}} & {in_wt_data79, in_wt_data78});
    in_wt_data_int16_38 = ({16{cfg_is_int16_d1[38]}} & {in_wt_data77, in_wt_data76});
    in_wt_data_int16_37 = ({16{cfg_is_int16_d1[37]}} & {in_wt_data75, in_wt_data74});
    in_wt_data_int16_36 = ({16{cfg_is_int16_d1[36]}} & {in_wt_data73, in_wt_data72});
    in_wt_data_int16_35 = ({16{cfg_is_int16_d1[35]}} & {in_wt_data71, in_wt_data70});
    in_wt_data_int16_34 = ({16{cfg_is_int16_d1[34]}} & {in_wt_data69, in_wt_data68});
    in_wt_data_int16_33 = ({16{cfg_is_int16_d1[33]}} & {in_wt_data67, in_wt_data66});
    in_wt_data_int16_32 = ({16{cfg_is_int16_d1[32]}} & {in_wt_data65, in_wt_data64});
    in_wt_data_int16_31 = ({16{cfg_is_int16_d1[31]}} & {in_wt_data63, in_wt_data62});
    in_wt_data_int16_30 = ({16{cfg_is_int16_d1[30]}} & {in_wt_data61, in_wt_data60});
    in_wt_data_int16_29 = ({16{cfg_is_int16_d1[29]}} & {in_wt_data59, in_wt_data58});
    in_wt_data_int16_28 = ({16{cfg_is_int16_d1[28]}} & {in_wt_data57, in_wt_data56});
    in_wt_data_int16_27 = ({16{cfg_is_int16_d1[27]}} & {in_wt_data55, in_wt_data54});
    in_wt_data_int16_26 = ({16{cfg_is_int16_d1[26]}} & {in_wt_data53, in_wt_data52});
    in_wt_data_int16_25 = ({16{cfg_is_int16_d1[25]}} & {in_wt_data51, in_wt_data50});
    in_wt_data_int16_24 = ({16{cfg_is_int16_d1[24]}} & {in_wt_data49, in_wt_data48});
    in_wt_data_int16_23 = ({16{cfg_is_int16_d1[23]}} & {in_wt_data47, in_wt_data46});
    in_wt_data_int16_22 = ({16{cfg_is_int16_d1[22]}} & {in_wt_data45, in_wt_data44});
    in_wt_data_int16_21 = ({16{cfg_is_int16_d1[21]}} & {in_wt_data43, in_wt_data42});
    in_wt_data_int16_20 = ({16{cfg_is_int16_d1[20]}} & {in_wt_data41, in_wt_data40});
    in_wt_data_int16_19 = ({16{cfg_is_int16_d1[19]}} & {in_wt_data39, in_wt_data38});
    in_wt_data_int16_18 = ({16{cfg_is_int16_d1[18]}} & {in_wt_data37, in_wt_data36});
    in_wt_data_int16_17 = ({16{cfg_is_int16_d1[17]}} & {in_wt_data35, in_wt_data34});
    in_wt_data_int16_16 = ({16{cfg_is_int16_d1[16]}} & {in_wt_data33, in_wt_data32});
    in_wt_data_int16_15 = ({16{cfg_is_int16_d1[15]}} & {in_wt_data31, in_wt_data30});
    in_wt_data_int16_14 = ({16{cfg_is_int16_d1[14]}} & {in_wt_data29, in_wt_data28});
    in_wt_data_int16_13 = ({16{cfg_is_int16_d1[13]}} & {in_wt_data27, in_wt_data26});
    in_wt_data_int16_12 = ({16{cfg_is_int16_d1[12]}} & {in_wt_data25, in_wt_data24});
    in_wt_data_int16_11 = ({16{cfg_is_int16_d1[11]}} & {in_wt_data23, in_wt_data22});
    in_wt_data_int16_10 = ({16{cfg_is_int16_d1[10]}} & {in_wt_data21, in_wt_data20});
    in_wt_data_int16_9 = ({16{cfg_is_int16_d1[9]}} & {in_wt_data19, in_wt_data18});
    in_wt_data_int16_8 = ({16{cfg_is_int16_d1[8]}} & {in_wt_data17, in_wt_data16});
    in_wt_data_int16_7 = ({16{cfg_is_int16_d1[7]}} & {in_wt_data15, in_wt_data14});
    in_wt_data_int16_6 = ({16{cfg_is_int16_d1[6]}} & {in_wt_data13, in_wt_data12});
    in_wt_data_int16_5 = ({16{cfg_is_int16_d1[5]}} & {in_wt_data11, in_wt_data10});
    in_wt_data_int16_4 = ({16{cfg_is_int16_d1[4]}} & {in_wt_data9, in_wt_data8});
    in_wt_data_int16_3 = ({16{cfg_is_int16_d1[3]}} & {in_wt_data7, in_wt_data6});
    in_wt_data_int16_2 = ({16{cfg_is_int16_d1[2]}} & {in_wt_data5, in_wt_data4});
    in_wt_data_int16_1 = ({16{cfg_is_int16_d1[1]}} & {in_wt_data3, in_wt_data2});
    in_wt_data_int16_0 = ({16{cfg_is_int16_d1[0]}} & {in_wt_data1, in_wt_data0});
end



always @(
  in_wt_data_int16_63
  or in_wt_data_int16_62
  or in_wt_data_int16_61
  or in_wt_data_int16_60
  or in_wt_data_int16_59
  or in_wt_data_int16_58
  or in_wt_data_int16_57
  or in_wt_data_int16_56
  or in_wt_data_int16_55
  or in_wt_data_int16_54
  or in_wt_data_int16_53
  or in_wt_data_int16_52
  or in_wt_data_int16_51
  or in_wt_data_int16_50
  or in_wt_data_int16_49
  or in_wt_data_int16_48
  or in_wt_data_int16_47
  or in_wt_data_int16_46
  or in_wt_data_int16_45
  or in_wt_data_int16_44
  or in_wt_data_int16_43
  or in_wt_data_int16_42
  or in_wt_data_int16_41
  or in_wt_data_int16_40
  or in_wt_data_int16_39
  or in_wt_data_int16_38
  or in_wt_data_int16_37
  or in_wt_data_int16_36
  or in_wt_data_int16_35
  or in_wt_data_int16_34
  or in_wt_data_int16_33
  or in_wt_data_int16_32
  or in_wt_data_int16_31
  or in_wt_data_int16_30
  or in_wt_data_int16_29
  or in_wt_data_int16_28
  or in_wt_data_int16_27
  or in_wt_data_int16_26
  or in_wt_data_int16_25
  or in_wt_data_int16_24
  or in_wt_data_int16_23
  or in_wt_data_int16_22
  or in_wt_data_int16_21
  or in_wt_data_int16_20
  or in_wt_data_int16_19
  or in_wt_data_int16_18
  or in_wt_data_int16_17
  or in_wt_data_int16_16
  or in_wt_data_int16_15
  or in_wt_data_int16_14
  or in_wt_data_int16_13
  or in_wt_data_int16_12
  or in_wt_data_int16_11
  or in_wt_data_int16_10
  or in_wt_data_int16_9
  or in_wt_data_int16_8
  or in_wt_data_int16_7
  or in_wt_data_int16_6
  or in_wt_data_int16_5
  or in_wt_data_int16_4
  or in_wt_data_int16_3
  or in_wt_data_int16_2
  or in_wt_data_int16_1
  or in_wt_data_int16_0
  ) begin
    in_wt_data_int16 = {in_wt_data_int16_63, in_wt_data_int16_62, in_wt_data_int16_61, in_wt_data_int16_60, in_wt_data_int16_59, in_wt_data_int16_58, in_wt_data_int16_57, in_wt_data_int16_56, in_wt_data_int16_55, in_wt_data_int16_54, in_wt_data_int16_53, in_wt_data_int16_52, in_wt_data_int16_51, in_wt_data_int16_50, in_wt_data_int16_49, in_wt_data_int16_48, in_wt_data_int16_47, in_wt_data_int16_46, in_wt_data_int16_45, in_wt_data_int16_44, in_wt_data_int16_43, in_wt_data_int16_42, in_wt_data_int16_41, in_wt_data_int16_40, in_wt_data_int16_39, in_wt_data_int16_38, in_wt_data_int16_37, in_wt_data_int16_36, in_wt_data_int16_35, in_wt_data_int16_34, in_wt_data_int16_33, in_wt_data_int16_32, in_wt_data_int16_31, in_wt_data_int16_30, in_wt_data_int16_29, in_wt_data_int16_28, in_wt_data_int16_27, in_wt_data_int16_26, in_wt_data_int16_25, in_wt_data_int16_24, in_wt_data_int16_23, in_wt_data_int16_22, in_wt_data_int16_21, in_wt_data_int16_20, in_wt_data_int16_19, in_wt_data_int16_18, in_wt_data_int16_17, in_wt_data_int16_16, in_wt_data_int16_15, in_wt_data_int16_14, in_wt_data_int16_13, in_wt_data_int16_12, in_wt_data_int16_11, in_wt_data_int16_10, in_wt_data_int16_9, in_wt_data_int16_8, in_wt_data_int16_7, in_wt_data_int16_6, in_wt_data_int16_5, in_wt_data_int16_4, in_wt_data_int16_3, in_wt_data_int16_2, in_wt_data_int16_1, in_wt_data_int16_0};
end

//////////////// in_wt_data_int8 ////////////////
always @(
  cfg_is_int8_d1
  or in_wt_data127
  or in_wt_data63
  or in_wt_data126
  or in_wt_data62
  or in_wt_data125
  or in_wt_data61
  or in_wt_data124
  or in_wt_data60
  or in_wt_data123
  or in_wt_data59
  or in_wt_data122
  or in_wt_data58
  or in_wt_data121
  or in_wt_data57
  or in_wt_data120
  or in_wt_data56
  or in_wt_data119
  or in_wt_data55
  or in_wt_data118
  or in_wt_data54
  or in_wt_data117
  or in_wt_data53
  or in_wt_data116
  or in_wt_data52
  or in_wt_data115
  or in_wt_data51
  or in_wt_data114
  or in_wt_data50
  or in_wt_data113
  or in_wt_data49
  or in_wt_data112
  or in_wt_data48
  or in_wt_data111
  or in_wt_data47
  or in_wt_data110
  or in_wt_data46
  or in_wt_data109
  or in_wt_data45
  or in_wt_data108
  or in_wt_data44
  or in_wt_data107
  or in_wt_data43
  or in_wt_data106
  or in_wt_data42
  or in_wt_data105
  or in_wt_data41
  or in_wt_data104
  or in_wt_data40
  or in_wt_data103
  or in_wt_data39
  or in_wt_data102
  or in_wt_data38
  or in_wt_data101
  or in_wt_data37
  or in_wt_data100
  or in_wt_data36
  or in_wt_data99
  or in_wt_data35
  or in_wt_data98
  or in_wt_data34
  or in_wt_data97
  or in_wt_data33
  or in_wt_data96
  or in_wt_data32
  or in_wt_data95
  or in_wt_data31
  or in_wt_data94
  or in_wt_data30
  or in_wt_data93
  or in_wt_data29
  or in_wt_data92
  or in_wt_data28
  or in_wt_data91
  or in_wt_data27
  or in_wt_data90
  or in_wt_data26
  or in_wt_data89
  or in_wt_data25
  or in_wt_data88
  or in_wt_data24
  or in_wt_data87
  or in_wt_data23
  or in_wt_data86
  or in_wt_data22
  or in_wt_data85
  or in_wt_data21
  or in_wt_data84
  or in_wt_data20
  or in_wt_data83
  or in_wt_data19
  or in_wt_data82
  or in_wt_data18
  or in_wt_data81
  or in_wt_data17
  or in_wt_data80
  or in_wt_data16
  or in_wt_data79
  or in_wt_data15
  or in_wt_data78
  or in_wt_data14
  or in_wt_data77
  or in_wt_data13
  or in_wt_data76
  or in_wt_data12
  or in_wt_data75
  or in_wt_data11
  or in_wt_data74
  or in_wt_data10
  or in_wt_data73
  or in_wt_data9
  or in_wt_data72
  or in_wt_data8
  or in_wt_data71
  or in_wt_data7
  or in_wt_data70
  or in_wt_data6
  or in_wt_data69
  or in_wt_data5
  or in_wt_data68
  or in_wt_data4
  or in_wt_data67
  or in_wt_data3
  or in_wt_data66
  or in_wt_data2
  or in_wt_data65
  or in_wt_data1
  or in_wt_data64
  or in_wt_data0
  ) begin
    in_wt_data_int8_63 = ({16{cfg_is_int8_d1[63]}} & {in_wt_data127, in_wt_data63});
    in_wt_data_int8_62 = ({16{cfg_is_int8_d1[62]}} & {in_wt_data126, in_wt_data62});
    in_wt_data_int8_61 = ({16{cfg_is_int8_d1[61]}} & {in_wt_data125, in_wt_data61});
    in_wt_data_int8_60 = ({16{cfg_is_int8_d1[60]}} & {in_wt_data124, in_wt_data60});
    in_wt_data_int8_59 = ({16{cfg_is_int8_d1[59]}} & {in_wt_data123, in_wt_data59});
    in_wt_data_int8_58 = ({16{cfg_is_int8_d1[58]}} & {in_wt_data122, in_wt_data58});
    in_wt_data_int8_57 = ({16{cfg_is_int8_d1[57]}} & {in_wt_data121, in_wt_data57});
    in_wt_data_int8_56 = ({16{cfg_is_int8_d1[56]}} & {in_wt_data120, in_wt_data56});
    in_wt_data_int8_55 = ({16{cfg_is_int8_d1[55]}} & {in_wt_data119, in_wt_data55});
    in_wt_data_int8_54 = ({16{cfg_is_int8_d1[54]}} & {in_wt_data118, in_wt_data54});
    in_wt_data_int8_53 = ({16{cfg_is_int8_d1[53]}} & {in_wt_data117, in_wt_data53});
    in_wt_data_int8_52 = ({16{cfg_is_int8_d1[52]}} & {in_wt_data116, in_wt_data52});
    in_wt_data_int8_51 = ({16{cfg_is_int8_d1[51]}} & {in_wt_data115, in_wt_data51});
    in_wt_data_int8_50 = ({16{cfg_is_int8_d1[50]}} & {in_wt_data114, in_wt_data50});
    in_wt_data_int8_49 = ({16{cfg_is_int8_d1[49]}} & {in_wt_data113, in_wt_data49});
    in_wt_data_int8_48 = ({16{cfg_is_int8_d1[48]}} & {in_wt_data112, in_wt_data48});
    in_wt_data_int8_47 = ({16{cfg_is_int8_d1[47]}} & {in_wt_data111, in_wt_data47});
    in_wt_data_int8_46 = ({16{cfg_is_int8_d1[46]}} & {in_wt_data110, in_wt_data46});
    in_wt_data_int8_45 = ({16{cfg_is_int8_d1[45]}} & {in_wt_data109, in_wt_data45});
    in_wt_data_int8_44 = ({16{cfg_is_int8_d1[44]}} & {in_wt_data108, in_wt_data44});
    in_wt_data_int8_43 = ({16{cfg_is_int8_d1[43]}} & {in_wt_data107, in_wt_data43});
    in_wt_data_int8_42 = ({16{cfg_is_int8_d1[42]}} & {in_wt_data106, in_wt_data42});
    in_wt_data_int8_41 = ({16{cfg_is_int8_d1[41]}} & {in_wt_data105, in_wt_data41});
    in_wt_data_int8_40 = ({16{cfg_is_int8_d1[40]}} & {in_wt_data104, in_wt_data40});
    in_wt_data_int8_39 = ({16{cfg_is_int8_d1[39]}} & {in_wt_data103, in_wt_data39});
    in_wt_data_int8_38 = ({16{cfg_is_int8_d1[38]}} & {in_wt_data102, in_wt_data38});
    in_wt_data_int8_37 = ({16{cfg_is_int8_d1[37]}} & {in_wt_data101, in_wt_data37});
    in_wt_data_int8_36 = ({16{cfg_is_int8_d1[36]}} & {in_wt_data100, in_wt_data36});
    in_wt_data_int8_35 = ({16{cfg_is_int8_d1[35]}} & {in_wt_data99, in_wt_data35});
    in_wt_data_int8_34 = ({16{cfg_is_int8_d1[34]}} & {in_wt_data98, in_wt_data34});
    in_wt_data_int8_33 = ({16{cfg_is_int8_d1[33]}} & {in_wt_data97, in_wt_data33});
    in_wt_data_int8_32 = ({16{cfg_is_int8_d1[32]}} & {in_wt_data96, in_wt_data32});
    in_wt_data_int8_31 = ({16{cfg_is_int8_d1[31]}} & {in_wt_data95, in_wt_data31});
    in_wt_data_int8_30 = ({16{cfg_is_int8_d1[30]}} & {in_wt_data94, in_wt_data30});
    in_wt_data_int8_29 = ({16{cfg_is_int8_d1[29]}} & {in_wt_data93, in_wt_data29});
    in_wt_data_int8_28 = ({16{cfg_is_int8_d1[28]}} & {in_wt_data92, in_wt_data28});
    in_wt_data_int8_27 = ({16{cfg_is_int8_d1[27]}} & {in_wt_data91, in_wt_data27});
    in_wt_data_int8_26 = ({16{cfg_is_int8_d1[26]}} & {in_wt_data90, in_wt_data26});
    in_wt_data_int8_25 = ({16{cfg_is_int8_d1[25]}} & {in_wt_data89, in_wt_data25});
    in_wt_data_int8_24 = ({16{cfg_is_int8_d1[24]}} & {in_wt_data88, in_wt_data24});
    in_wt_data_int8_23 = ({16{cfg_is_int8_d1[23]}} & {in_wt_data87, in_wt_data23});
    in_wt_data_int8_22 = ({16{cfg_is_int8_d1[22]}} & {in_wt_data86, in_wt_data22});
    in_wt_data_int8_21 = ({16{cfg_is_int8_d1[21]}} & {in_wt_data85, in_wt_data21});
    in_wt_data_int8_20 = ({16{cfg_is_int8_d1[20]}} & {in_wt_data84, in_wt_data20});
    in_wt_data_int8_19 = ({16{cfg_is_int8_d1[19]}} & {in_wt_data83, in_wt_data19});
    in_wt_data_int8_18 = ({16{cfg_is_int8_d1[18]}} & {in_wt_data82, in_wt_data18});
    in_wt_data_int8_17 = ({16{cfg_is_int8_d1[17]}} & {in_wt_data81, in_wt_data17});
    in_wt_data_int8_16 = ({16{cfg_is_int8_d1[16]}} & {in_wt_data80, in_wt_data16});
    in_wt_data_int8_15 = ({16{cfg_is_int8_d1[15]}} & {in_wt_data79, in_wt_data15});
    in_wt_data_int8_14 = ({16{cfg_is_int8_d1[14]}} & {in_wt_data78, in_wt_data14});
    in_wt_data_int8_13 = ({16{cfg_is_int8_d1[13]}} & {in_wt_data77, in_wt_data13});
    in_wt_data_int8_12 = ({16{cfg_is_int8_d1[12]}} & {in_wt_data76, in_wt_data12});
    in_wt_data_int8_11 = ({16{cfg_is_int8_d1[11]}} & {in_wt_data75, in_wt_data11});
    in_wt_data_int8_10 = ({16{cfg_is_int8_d1[10]}} & {in_wt_data74, in_wt_data10});
    in_wt_data_int8_9 = ({16{cfg_is_int8_d1[9]}} & {in_wt_data73, in_wt_data9});
    in_wt_data_int8_8 = ({16{cfg_is_int8_d1[8]}} & {in_wt_data72, in_wt_data8});
    in_wt_data_int8_7 = ({16{cfg_is_int8_d1[7]}} & {in_wt_data71, in_wt_data7});
    in_wt_data_int8_6 = ({16{cfg_is_int8_d1[6]}} & {in_wt_data70, in_wt_data6});
    in_wt_data_int8_5 = ({16{cfg_is_int8_d1[5]}} & {in_wt_data69, in_wt_data5});
    in_wt_data_int8_4 = ({16{cfg_is_int8_d1[4]}} & {in_wt_data68, in_wt_data4});
    in_wt_data_int8_3 = ({16{cfg_is_int8_d1[3]}} & {in_wt_data67, in_wt_data3});
    in_wt_data_int8_2 = ({16{cfg_is_int8_d1[2]}} & {in_wt_data66, in_wt_data2});
    in_wt_data_int8_1 = ({16{cfg_is_int8_d1[1]}} & {in_wt_data65, in_wt_data1});
    in_wt_data_int8_0 = ({16{cfg_is_int8_d1[0]}} & {in_wt_data64, in_wt_data0});
end


always @(
  in_wt_mask
  ) begin
    in_wt_mask_int8 = {in_wt_mask[127], in_wt_mask[63], in_wt_mask[126], in_wt_mask[62], in_wt_mask[125], in_wt_mask[61], in_wt_mask[124], in_wt_mask[60], in_wt_mask[123], in_wt_mask[59], in_wt_mask[122], in_wt_mask[58], in_wt_mask[121], in_wt_mask[57], in_wt_mask[120], in_wt_mask[56],
                       in_wt_mask[119], in_wt_mask[55], in_wt_mask[118], in_wt_mask[54], in_wt_mask[117], in_wt_mask[53], in_wt_mask[116], in_wt_mask[52], in_wt_mask[115], in_wt_mask[51], in_wt_mask[114], in_wt_mask[50], in_wt_mask[113], in_wt_mask[49], in_wt_mask[112], in_wt_mask[48],
                       in_wt_mask[111], in_wt_mask[47], in_wt_mask[110], in_wt_mask[46], in_wt_mask[109], in_wt_mask[45], in_wt_mask[108], in_wt_mask[44], in_wt_mask[107], in_wt_mask[43], in_wt_mask[106], in_wt_mask[42], in_wt_mask[105], in_wt_mask[41], in_wt_mask[104], in_wt_mask[40],
                       in_wt_mask[103], in_wt_mask[39], in_wt_mask[102], in_wt_mask[38], in_wt_mask[101], in_wt_mask[37], in_wt_mask[100], in_wt_mask[36], in_wt_mask[99], in_wt_mask[35], in_wt_mask[98], in_wt_mask[34], in_wt_mask[97], in_wt_mask[33], in_wt_mask[96], in_wt_mask[32],
                       in_wt_mask[95], in_wt_mask[31], in_wt_mask[94], in_wt_mask[30], in_wt_mask[93], in_wt_mask[29], in_wt_mask[92], in_wt_mask[28], in_wt_mask[91], in_wt_mask[27], in_wt_mask[90], in_wt_mask[26], in_wt_mask[89], in_wt_mask[25], in_wt_mask[88], in_wt_mask[24],
                       in_wt_mask[87], in_wt_mask[23], in_wt_mask[86], in_wt_mask[22], in_wt_mask[85], in_wt_mask[21], in_wt_mask[84], in_wt_mask[20], in_wt_mask[83], in_wt_mask[19], in_wt_mask[82], in_wt_mask[18], in_wt_mask[81], in_wt_mask[17], in_wt_mask[80], in_wt_mask[16],
                       in_wt_mask[79], in_wt_mask[15], in_wt_mask[78], in_wt_mask[14], in_wt_mask[77], in_wt_mask[13], in_wt_mask[76], in_wt_mask[12], in_wt_mask[75], in_wt_mask[11], in_wt_mask[74], in_wt_mask[10], in_wt_mask[73], in_wt_mask[9], in_wt_mask[72], in_wt_mask[8],
                       in_wt_mask[71], in_wt_mask[7], in_wt_mask[70], in_wt_mask[6], in_wt_mask[69], in_wt_mask[5], in_wt_mask[68], in_wt_mask[4], in_wt_mask[67], in_wt_mask[3], in_wt_mask[66], in_wt_mask[2], in_wt_mask[65], in_wt_mask[1], in_wt_mask[64], in_wt_mask[0]};
end



always @(
  in_wt_data_int8_63
  or in_wt_data_int8_62
  or in_wt_data_int8_61
  or in_wt_data_int8_60
  or in_wt_data_int8_59
  or in_wt_data_int8_58
  or in_wt_data_int8_57
  or in_wt_data_int8_56
  or in_wt_data_int8_55
  or in_wt_data_int8_54
  or in_wt_data_int8_53
  or in_wt_data_int8_52
  or in_wt_data_int8_51
  or in_wt_data_int8_50
  or in_wt_data_int8_49
  or in_wt_data_int8_48
  or in_wt_data_int8_47
  or in_wt_data_int8_46
  or in_wt_data_int8_45
  or in_wt_data_int8_44
  or in_wt_data_int8_43
  or in_wt_data_int8_42
  or in_wt_data_int8_41
  or in_wt_data_int8_40
  or in_wt_data_int8_39
  or in_wt_data_int8_38
  or in_wt_data_int8_37
  or in_wt_data_int8_36
  or in_wt_data_int8_35
  or in_wt_data_int8_34
  or in_wt_data_int8_33
  or in_wt_data_int8_32
  or in_wt_data_int8_31
  or in_wt_data_int8_30
  or in_wt_data_int8_29
  or in_wt_data_int8_28
  or in_wt_data_int8_27
  or in_wt_data_int8_26
  or in_wt_data_int8_25
  or in_wt_data_int8_24
  or in_wt_data_int8_23
  or in_wt_data_int8_22
  or in_wt_data_int8_21
  or in_wt_data_int8_20
  or in_wt_data_int8_19
  or in_wt_data_int8_18
  or in_wt_data_int8_17
  or in_wt_data_int8_16
  or in_wt_data_int8_15
  or in_wt_data_int8_14
  or in_wt_data_int8_13
  or in_wt_data_int8_12
  or in_wt_data_int8_11
  or in_wt_data_int8_10
  or in_wt_data_int8_9
  or in_wt_data_int8_8
  or in_wt_data_int8_7
  or in_wt_data_int8_6
  or in_wt_data_int8_5
  or in_wt_data_int8_4
  or in_wt_data_int8_3
  or in_wt_data_int8_2
  or in_wt_data_int8_1
  or in_wt_data_int8_0
  ) begin
    in_wt_data_int8 = {in_wt_data_int8_63, in_wt_data_int8_62, in_wt_data_int8_61, in_wt_data_int8_60, in_wt_data_int8_59, in_wt_data_int8_58, in_wt_data_int8_57, in_wt_data_int8_56, in_wt_data_int8_55, in_wt_data_int8_54, in_wt_data_int8_53, in_wt_data_int8_52, in_wt_data_int8_51, in_wt_data_int8_50, in_wt_data_int8_49, in_wt_data_int8_48, in_wt_data_int8_47, in_wt_data_int8_46, in_wt_data_int8_45, in_wt_data_int8_44, in_wt_data_int8_43, in_wt_data_int8_42, in_wt_data_int8_41, in_wt_data_int8_40, in_wt_data_int8_39, in_wt_data_int8_38, in_wt_data_int8_37, in_wt_data_int8_36, in_wt_data_int8_35, in_wt_data_int8_34, in_wt_data_int8_33, in_wt_data_int8_32, in_wt_data_int8_31, in_wt_data_int8_30, in_wt_data_int8_29, in_wt_data_int8_28, in_wt_data_int8_27, in_wt_data_int8_26, in_wt_data_int8_25, in_wt_data_int8_24, in_wt_data_int8_23, in_wt_data_int8_22, in_wt_data_int8_21, in_wt_data_int8_20, in_wt_data_int8_19, in_wt_data_int8_18, in_wt_data_int8_17, in_wt_data_int8_16, in_wt_data_int8_15, in_wt_data_int8_14, in_wt_data_int8_13, in_wt_data_int8_12, in_wt_data_int8_11, in_wt_data_int8_10, in_wt_data_int8_9, in_wt_data_int8_8, in_wt_data_int8_7, in_wt_data_int8_6, in_wt_data_int8_5, in_wt_data_int8_4, in_wt_data_int8_3, in_wt_data_int8_2, in_wt_data_int8_1, in_wt_data_int8_0};
end

//////////////// in_wt_data_fp16 ////////////////
always @(
  cfg_is_fp16_d1
  or in_wt_data_pack
  or in_wt_mask
  ) begin
    in_wt_nan[63] = cfg_is_fp16_d1[63] & (&in_wt_data_pack[1022:1018]) & (|in_wt_data_pack[1017:1008]) & in_wt_mask[126];
    in_wt_nan[62] = cfg_is_fp16_d1[62] & (&in_wt_data_pack[1006:1002]) & (|in_wt_data_pack[1001:992]) & in_wt_mask[124];
    in_wt_nan[61] = cfg_is_fp16_d1[61] & (&in_wt_data_pack[990:986]) & (|in_wt_data_pack[985:976]) & in_wt_mask[122];
    in_wt_nan[60] = cfg_is_fp16_d1[60] & (&in_wt_data_pack[974:970]) & (|in_wt_data_pack[969:960]) & in_wt_mask[120];
    in_wt_nan[59] = cfg_is_fp16_d1[59] & (&in_wt_data_pack[958:954]) & (|in_wt_data_pack[953:944]) & in_wt_mask[118];
    in_wt_nan[58] = cfg_is_fp16_d1[58] & (&in_wt_data_pack[942:938]) & (|in_wt_data_pack[937:928]) & in_wt_mask[116];
    in_wt_nan[57] = cfg_is_fp16_d1[57] & (&in_wt_data_pack[926:922]) & (|in_wt_data_pack[921:912]) & in_wt_mask[114];
    in_wt_nan[56] = cfg_is_fp16_d1[56] & (&in_wt_data_pack[910:906]) & (|in_wt_data_pack[905:896]) & in_wt_mask[112];
    in_wt_nan[55] = cfg_is_fp16_d1[55] & (&in_wt_data_pack[894:890]) & (|in_wt_data_pack[889:880]) & in_wt_mask[110];
    in_wt_nan[54] = cfg_is_fp16_d1[54] & (&in_wt_data_pack[878:874]) & (|in_wt_data_pack[873:864]) & in_wt_mask[108];
    in_wt_nan[53] = cfg_is_fp16_d1[53] & (&in_wt_data_pack[862:858]) & (|in_wt_data_pack[857:848]) & in_wt_mask[106];
    in_wt_nan[52] = cfg_is_fp16_d1[52] & (&in_wt_data_pack[846:842]) & (|in_wt_data_pack[841:832]) & in_wt_mask[104];
    in_wt_nan[51] = cfg_is_fp16_d1[51] & (&in_wt_data_pack[830:826]) & (|in_wt_data_pack[825:816]) & in_wt_mask[102];
    in_wt_nan[50] = cfg_is_fp16_d1[50] & (&in_wt_data_pack[814:810]) & (|in_wt_data_pack[809:800]) & in_wt_mask[100];
    in_wt_nan[49] = cfg_is_fp16_d1[49] & (&in_wt_data_pack[798:794]) & (|in_wt_data_pack[793:784]) & in_wt_mask[98];
    in_wt_nan[48] = cfg_is_fp16_d1[48] & (&in_wt_data_pack[782:778]) & (|in_wt_data_pack[777:768]) & in_wt_mask[96];
    in_wt_nan[47] = cfg_is_fp16_d1[47] & (&in_wt_data_pack[766:762]) & (|in_wt_data_pack[761:752]) & in_wt_mask[94];
    in_wt_nan[46] = cfg_is_fp16_d1[46] & (&in_wt_data_pack[750:746]) & (|in_wt_data_pack[745:736]) & in_wt_mask[92];
    in_wt_nan[45] = cfg_is_fp16_d1[45] & (&in_wt_data_pack[734:730]) & (|in_wt_data_pack[729:720]) & in_wt_mask[90];
    in_wt_nan[44] = cfg_is_fp16_d1[44] & (&in_wt_data_pack[718:714]) & (|in_wt_data_pack[713:704]) & in_wt_mask[88];
    in_wt_nan[43] = cfg_is_fp16_d1[43] & (&in_wt_data_pack[702:698]) & (|in_wt_data_pack[697:688]) & in_wt_mask[86];
    in_wt_nan[42] = cfg_is_fp16_d1[42] & (&in_wt_data_pack[686:682]) & (|in_wt_data_pack[681:672]) & in_wt_mask[84];
    in_wt_nan[41] = cfg_is_fp16_d1[41] & (&in_wt_data_pack[670:666]) & (|in_wt_data_pack[665:656]) & in_wt_mask[82];
    in_wt_nan[40] = cfg_is_fp16_d1[40] & (&in_wt_data_pack[654:650]) & (|in_wt_data_pack[649:640]) & in_wt_mask[80];
    in_wt_nan[39] = cfg_is_fp16_d1[39] & (&in_wt_data_pack[638:634]) & (|in_wt_data_pack[633:624]) & in_wt_mask[78];
    in_wt_nan[38] = cfg_is_fp16_d1[38] & (&in_wt_data_pack[622:618]) & (|in_wt_data_pack[617:608]) & in_wt_mask[76];
    in_wt_nan[37] = cfg_is_fp16_d1[37] & (&in_wt_data_pack[606:602]) & (|in_wt_data_pack[601:592]) & in_wt_mask[74];
    in_wt_nan[36] = cfg_is_fp16_d1[36] & (&in_wt_data_pack[590:586]) & (|in_wt_data_pack[585:576]) & in_wt_mask[72];
    in_wt_nan[35] = cfg_is_fp16_d1[35] & (&in_wt_data_pack[574:570]) & (|in_wt_data_pack[569:560]) & in_wt_mask[70];
    in_wt_nan[34] = cfg_is_fp16_d1[34] & (&in_wt_data_pack[558:554]) & (|in_wt_data_pack[553:544]) & in_wt_mask[68];
    in_wt_nan[33] = cfg_is_fp16_d1[33] & (&in_wt_data_pack[542:538]) & (|in_wt_data_pack[537:528]) & in_wt_mask[66];
    in_wt_nan[32] = cfg_is_fp16_d1[32] & (&in_wt_data_pack[526:522]) & (|in_wt_data_pack[521:512]) & in_wt_mask[64];
    in_wt_nan[31] = cfg_is_fp16_d1[31] & (&in_wt_data_pack[510:506]) & (|in_wt_data_pack[505:496]) & in_wt_mask[62];
    in_wt_nan[30] = cfg_is_fp16_d1[30] & (&in_wt_data_pack[494:490]) & (|in_wt_data_pack[489:480]) & in_wt_mask[60];
    in_wt_nan[29] = cfg_is_fp16_d1[29] & (&in_wt_data_pack[478:474]) & (|in_wt_data_pack[473:464]) & in_wt_mask[58];
    in_wt_nan[28] = cfg_is_fp16_d1[28] & (&in_wt_data_pack[462:458]) & (|in_wt_data_pack[457:448]) & in_wt_mask[56];
    in_wt_nan[27] = cfg_is_fp16_d1[27] & (&in_wt_data_pack[446:442]) & (|in_wt_data_pack[441:432]) & in_wt_mask[54];
    in_wt_nan[26] = cfg_is_fp16_d1[26] & (&in_wt_data_pack[430:426]) & (|in_wt_data_pack[425:416]) & in_wt_mask[52];
    in_wt_nan[25] = cfg_is_fp16_d1[25] & (&in_wt_data_pack[414:410]) & (|in_wt_data_pack[409:400]) & in_wt_mask[50];
    in_wt_nan[24] = cfg_is_fp16_d1[24] & (&in_wt_data_pack[398:394]) & (|in_wt_data_pack[393:384]) & in_wt_mask[48];
    in_wt_nan[23] = cfg_is_fp16_d1[23] & (&in_wt_data_pack[382:378]) & (|in_wt_data_pack[377:368]) & in_wt_mask[46];
    in_wt_nan[22] = cfg_is_fp16_d1[22] & (&in_wt_data_pack[366:362]) & (|in_wt_data_pack[361:352]) & in_wt_mask[44];
    in_wt_nan[21] = cfg_is_fp16_d1[21] & (&in_wt_data_pack[350:346]) & (|in_wt_data_pack[345:336]) & in_wt_mask[42];
    in_wt_nan[20] = cfg_is_fp16_d1[20] & (&in_wt_data_pack[334:330]) & (|in_wt_data_pack[329:320]) & in_wt_mask[40];
    in_wt_nan[19] = cfg_is_fp16_d1[19] & (&in_wt_data_pack[318:314]) & (|in_wt_data_pack[313:304]) & in_wt_mask[38];
    in_wt_nan[18] = cfg_is_fp16_d1[18] & (&in_wt_data_pack[302:298]) & (|in_wt_data_pack[297:288]) & in_wt_mask[36];
    in_wt_nan[17] = cfg_is_fp16_d1[17] & (&in_wt_data_pack[286:282]) & (|in_wt_data_pack[281:272]) & in_wt_mask[34];
    in_wt_nan[16] = cfg_is_fp16_d1[16] & (&in_wt_data_pack[270:266]) & (|in_wt_data_pack[265:256]) & in_wt_mask[32];
    in_wt_nan[15] = cfg_is_fp16_d1[15] & (&in_wt_data_pack[254:250]) & (|in_wt_data_pack[249:240]) & in_wt_mask[30];
    in_wt_nan[14] = cfg_is_fp16_d1[14] & (&in_wt_data_pack[238:234]) & (|in_wt_data_pack[233:224]) & in_wt_mask[28];
    in_wt_nan[13] = cfg_is_fp16_d1[13] & (&in_wt_data_pack[222:218]) & (|in_wt_data_pack[217:208]) & in_wt_mask[26];
    in_wt_nan[12] = cfg_is_fp16_d1[12] & (&in_wt_data_pack[206:202]) & (|in_wt_data_pack[201:192]) & in_wt_mask[24];
    in_wt_nan[11] = cfg_is_fp16_d1[11] & (&in_wt_data_pack[190:186]) & (|in_wt_data_pack[185:176]) & in_wt_mask[22];
    in_wt_nan[10] = cfg_is_fp16_d1[10] & (&in_wt_data_pack[174:170]) & (|in_wt_data_pack[169:160]) & in_wt_mask[20];
    in_wt_nan[9] = cfg_is_fp16_d1[9] & (&in_wt_data_pack[158:154]) & (|in_wt_data_pack[153:144]) & in_wt_mask[18];
    in_wt_nan[8] = cfg_is_fp16_d1[8] & (&in_wt_data_pack[142:138]) & (|in_wt_data_pack[137:128]) & in_wt_mask[16];
    in_wt_nan[7] = cfg_is_fp16_d1[7] & (&in_wt_data_pack[126:122]) & (|in_wt_data_pack[121:112]) & in_wt_mask[14];
    in_wt_nan[6] = cfg_is_fp16_d1[6] & (&in_wt_data_pack[110:106]) & (|in_wt_data_pack[105:96]) & in_wt_mask[12];
    in_wt_nan[5] = cfg_is_fp16_d1[5] & (&in_wt_data_pack[94:90]) & (|in_wt_data_pack[89:80]) & in_wt_mask[10];
    in_wt_nan[4] = cfg_is_fp16_d1[4] & (&in_wt_data_pack[78:74]) & (|in_wt_data_pack[73:64]) & in_wt_mask[8];
    in_wt_nan[3] = cfg_is_fp16_d1[3] & (&in_wt_data_pack[62:58]) & (|in_wt_data_pack[57:48]) & in_wt_mask[6];
    in_wt_nan[2] = cfg_is_fp16_d1[2] & (&in_wt_data_pack[46:42]) & (|in_wt_data_pack[41:32]) & in_wt_mask[4];
    in_wt_nan[1] = cfg_is_fp16_d1[1] & (&in_wt_data_pack[30:26]) & (|in_wt_data_pack[25:16]) & in_wt_mask[2];
    in_wt_nan[0] = cfg_is_fp16_d1[0] & (&in_wt_data_pack[14:10]) & (|in_wt_data_pack[9:0]) & in_wt_mask[0];
end


always @(
  cfg_is_fp16_d1
  or in_wt_mask
  or in_wt_data_pack
  ) begin
    in_wt_exp[191:189] = {3{cfg_is_fp16_d1[63] & in_wt_mask[127]}} & (in_wt_data_pack[1022:1020]);
    in_wt_exp[188:186] = {3{cfg_is_fp16_d1[62] & in_wt_mask[125]}} & (in_wt_data_pack[1006:1004]);
    in_wt_exp[185:183] = {3{cfg_is_fp16_d1[61] & in_wt_mask[123]}} & (in_wt_data_pack[990:988]);
    in_wt_exp[182:180] = {3{cfg_is_fp16_d1[60] & in_wt_mask[121]}} & (in_wt_data_pack[974:972]);
    in_wt_exp[179:177] = {3{cfg_is_fp16_d1[59] & in_wt_mask[119]}} & (in_wt_data_pack[958:956]);
    in_wt_exp[176:174] = {3{cfg_is_fp16_d1[58] & in_wt_mask[117]}} & (in_wt_data_pack[942:940]);
    in_wt_exp[173:171] = {3{cfg_is_fp16_d1[57] & in_wt_mask[115]}} & (in_wt_data_pack[926:924]);
    in_wt_exp[170:168] = {3{cfg_is_fp16_d1[56] & in_wt_mask[113]}} & (in_wt_data_pack[910:908]);
    in_wt_exp[167:165] = {3{cfg_is_fp16_d1[55] & in_wt_mask[111]}} & (in_wt_data_pack[894:892]);
    in_wt_exp[164:162] = {3{cfg_is_fp16_d1[54] & in_wt_mask[109]}} & (in_wt_data_pack[878:876]);
    in_wt_exp[161:159] = {3{cfg_is_fp16_d1[53] & in_wt_mask[107]}} & (in_wt_data_pack[862:860]);
    in_wt_exp[158:156] = {3{cfg_is_fp16_d1[52] & in_wt_mask[105]}} & (in_wt_data_pack[846:844]);
    in_wt_exp[155:153] = {3{cfg_is_fp16_d1[51] & in_wt_mask[103]}} & (in_wt_data_pack[830:828]);
    in_wt_exp[152:150] = {3{cfg_is_fp16_d1[50] & in_wt_mask[101]}} & (in_wt_data_pack[814:812]);
    in_wt_exp[149:147] = {3{cfg_is_fp16_d1[49] & in_wt_mask[99]}} & (in_wt_data_pack[798:796]);
    in_wt_exp[146:144] = {3{cfg_is_fp16_d1[48] & in_wt_mask[97]}} & (in_wt_data_pack[782:780]);
    in_wt_exp[143:141] = {3{cfg_is_fp16_d1[47] & in_wt_mask[95]}} & (in_wt_data_pack[766:764]);
    in_wt_exp[140:138] = {3{cfg_is_fp16_d1[46] & in_wt_mask[93]}} & (in_wt_data_pack[750:748]);
    in_wt_exp[137:135] = {3{cfg_is_fp16_d1[45] & in_wt_mask[91]}} & (in_wt_data_pack[734:732]);
    in_wt_exp[134:132] = {3{cfg_is_fp16_d1[44] & in_wt_mask[89]}} & (in_wt_data_pack[718:716]);
    in_wt_exp[131:129] = {3{cfg_is_fp16_d1[43] & in_wt_mask[87]}} & (in_wt_data_pack[702:700]);
    in_wt_exp[128:126] = {3{cfg_is_fp16_d1[42] & in_wt_mask[85]}} & (in_wt_data_pack[686:684]);
    in_wt_exp[125:123] = {3{cfg_is_fp16_d1[41] & in_wt_mask[83]}} & (in_wt_data_pack[670:668]);
    in_wt_exp[122:120] = {3{cfg_is_fp16_d1[40] & in_wt_mask[81]}} & (in_wt_data_pack[654:652]);
    in_wt_exp[119:117] = {3{cfg_is_fp16_d1[39] & in_wt_mask[79]}} & (in_wt_data_pack[638:636]);
    in_wt_exp[116:114] = {3{cfg_is_fp16_d1[38] & in_wt_mask[77]}} & (in_wt_data_pack[622:620]);
    in_wt_exp[113:111] = {3{cfg_is_fp16_d1[37] & in_wt_mask[75]}} & (in_wt_data_pack[606:604]);
    in_wt_exp[110:108] = {3{cfg_is_fp16_d1[36] & in_wt_mask[73]}} & (in_wt_data_pack[590:588]);
    in_wt_exp[107:105] = {3{cfg_is_fp16_d1[35] & in_wt_mask[71]}} & (in_wt_data_pack[574:572]);
    in_wt_exp[104:102] = {3{cfg_is_fp16_d1[34] & in_wt_mask[69]}} & (in_wt_data_pack[558:556]);
    in_wt_exp[101:99] = {3{cfg_is_fp16_d1[33] & in_wt_mask[67]}} & (in_wt_data_pack[542:540]);
    in_wt_exp[98:96] = {3{cfg_is_fp16_d1[32] & in_wt_mask[65]}} & (in_wt_data_pack[526:524]);
    in_wt_exp[95:93] = {3{cfg_is_fp16_d1[31] & in_wt_mask[63]}} & (in_wt_data_pack[510:508]);
    in_wt_exp[92:90] = {3{cfg_is_fp16_d1[30] & in_wt_mask[61]}} & (in_wt_data_pack[494:492]);
    in_wt_exp[89:87] = {3{cfg_is_fp16_d1[29] & in_wt_mask[59]}} & (in_wt_data_pack[478:476]);
    in_wt_exp[86:84] = {3{cfg_is_fp16_d1[28] & in_wt_mask[57]}} & (in_wt_data_pack[462:460]);
    in_wt_exp[83:81] = {3{cfg_is_fp16_d1[27] & in_wt_mask[55]}} & (in_wt_data_pack[446:444]);
    in_wt_exp[80:78] = {3{cfg_is_fp16_d1[26] & in_wt_mask[53]}} & (in_wt_data_pack[430:428]);
    in_wt_exp[77:75] = {3{cfg_is_fp16_d1[25] & in_wt_mask[51]}} & (in_wt_data_pack[414:412]);
    in_wt_exp[74:72] = {3{cfg_is_fp16_d1[24] & in_wt_mask[49]}} & (in_wt_data_pack[398:396]);
    in_wt_exp[71:69] = {3{cfg_is_fp16_d1[23] & in_wt_mask[47]}} & (in_wt_data_pack[382:380]);
    in_wt_exp[68:66] = {3{cfg_is_fp16_d1[22] & in_wt_mask[45]}} & (in_wt_data_pack[366:364]);
    in_wt_exp[65:63] = {3{cfg_is_fp16_d1[21] & in_wt_mask[43]}} & (in_wt_data_pack[350:348]);
    in_wt_exp[62:60] = {3{cfg_is_fp16_d1[20] & in_wt_mask[41]}} & (in_wt_data_pack[334:332]);
    in_wt_exp[59:57] = {3{cfg_is_fp16_d1[19] & in_wt_mask[39]}} & (in_wt_data_pack[318:316]);
    in_wt_exp[56:54] = {3{cfg_is_fp16_d1[18] & in_wt_mask[37]}} & (in_wt_data_pack[302:300]);
    in_wt_exp[53:51] = {3{cfg_is_fp16_d1[17] & in_wt_mask[35]}} & (in_wt_data_pack[286:284]);
    in_wt_exp[50:48] = {3{cfg_is_fp16_d1[16] & in_wt_mask[33]}} & (in_wt_data_pack[270:268]);
    in_wt_exp[47:45] = {3{cfg_is_fp16_d1[15] & in_wt_mask[31]}} & (in_wt_data_pack[254:252]);
    in_wt_exp[44:42] = {3{cfg_is_fp16_d1[14] & in_wt_mask[29]}} & (in_wt_data_pack[238:236]);
    in_wt_exp[41:39] = {3{cfg_is_fp16_d1[13] & in_wt_mask[27]}} & (in_wt_data_pack[222:220]);
    in_wt_exp[38:36] = {3{cfg_is_fp16_d1[12] & in_wt_mask[25]}} & (in_wt_data_pack[206:204]);
    in_wt_exp[35:33] = {3{cfg_is_fp16_d1[11] & in_wt_mask[23]}} & (in_wt_data_pack[190:188]);
    in_wt_exp[32:30] = {3{cfg_is_fp16_d1[10] & in_wt_mask[21]}} & (in_wt_data_pack[174:172]);
    in_wt_exp[29:27] = {3{cfg_is_fp16_d1[9] & in_wt_mask[19]}} & (in_wt_data_pack[158:156]);
    in_wt_exp[26:24] = {3{cfg_is_fp16_d1[8] & in_wt_mask[17]}} & (in_wt_data_pack[142:140]);
    in_wt_exp[23:21] = {3{cfg_is_fp16_d1[7] & in_wt_mask[15]}} & (in_wt_data_pack[126:124]);
    in_wt_exp[20:18] = {3{cfg_is_fp16_d1[6] & in_wt_mask[13]}} & (in_wt_data_pack[110:108]);
    in_wt_exp[17:15] = {3{cfg_is_fp16_d1[5] & in_wt_mask[11]}} & (in_wt_data_pack[94:92]);
    in_wt_exp[14:12] = {3{cfg_is_fp16_d1[4] & in_wt_mask[9]}} & (in_wt_data_pack[78:76]);
    in_wt_exp[11:9] = {3{cfg_is_fp16_d1[3] & in_wt_mask[7]}} & (in_wt_data_pack[62:60]);
    in_wt_exp[8:6] = {3{cfg_is_fp16_d1[2] & in_wt_mask[5]}} & (in_wt_data_pack[46:44]);
    in_wt_exp[5:3] = {3{cfg_is_fp16_d1[1] & in_wt_mask[3]}} & (in_wt_data_pack[30:28]);
    in_wt_exp[2:0] = {3{cfg_is_fp16_d1[0] & in_wt_mask[1]}} & (in_wt_data_pack[14:12]);
end


always @(
  cfg_is_fp16_d1
  or in_wt_data_pack
  ) begin
    in_wt_norm[63] = cfg_is_fp16_d1[63] & (|in_wt_data_pack[1022:1018]);
    in_wt_norm[62] = cfg_is_fp16_d1[62] & (|in_wt_data_pack[1006:1002]);
    in_wt_norm[61] = cfg_is_fp16_d1[61] & (|in_wt_data_pack[990:986]);
    in_wt_norm[60] = cfg_is_fp16_d1[60] & (|in_wt_data_pack[974:970]);
    in_wt_norm[59] = cfg_is_fp16_d1[59] & (|in_wt_data_pack[958:954]);
    in_wt_norm[58] = cfg_is_fp16_d1[58] & (|in_wt_data_pack[942:938]);
    in_wt_norm[57] = cfg_is_fp16_d1[57] & (|in_wt_data_pack[926:922]);
    in_wt_norm[56] = cfg_is_fp16_d1[56] & (|in_wt_data_pack[910:906]);
    in_wt_norm[55] = cfg_is_fp16_d1[55] & (|in_wt_data_pack[894:890]);
    in_wt_norm[54] = cfg_is_fp16_d1[54] & (|in_wt_data_pack[878:874]);
    in_wt_norm[53] = cfg_is_fp16_d1[53] & (|in_wt_data_pack[862:858]);
    in_wt_norm[52] = cfg_is_fp16_d1[52] & (|in_wt_data_pack[846:842]);
    in_wt_norm[51] = cfg_is_fp16_d1[51] & (|in_wt_data_pack[830:826]);
    in_wt_norm[50] = cfg_is_fp16_d1[50] & (|in_wt_data_pack[814:810]);
    in_wt_norm[49] = cfg_is_fp16_d1[49] & (|in_wt_data_pack[798:794]);
    in_wt_norm[48] = cfg_is_fp16_d1[48] & (|in_wt_data_pack[782:778]);
    in_wt_norm[47] = cfg_is_fp16_d1[47] & (|in_wt_data_pack[766:762]);
    in_wt_norm[46] = cfg_is_fp16_d1[46] & (|in_wt_data_pack[750:746]);
    in_wt_norm[45] = cfg_is_fp16_d1[45] & (|in_wt_data_pack[734:730]);
    in_wt_norm[44] = cfg_is_fp16_d1[44] & (|in_wt_data_pack[718:714]);
    in_wt_norm[43] = cfg_is_fp16_d1[43] & (|in_wt_data_pack[702:698]);
    in_wt_norm[42] = cfg_is_fp16_d1[42] & (|in_wt_data_pack[686:682]);
    in_wt_norm[41] = cfg_is_fp16_d1[41] & (|in_wt_data_pack[670:666]);
    in_wt_norm[40] = cfg_is_fp16_d1[40] & (|in_wt_data_pack[654:650]);
    in_wt_norm[39] = cfg_is_fp16_d1[39] & (|in_wt_data_pack[638:634]);
    in_wt_norm[38] = cfg_is_fp16_d1[38] & (|in_wt_data_pack[622:618]);
    in_wt_norm[37] = cfg_is_fp16_d1[37] & (|in_wt_data_pack[606:602]);
    in_wt_norm[36] = cfg_is_fp16_d1[36] & (|in_wt_data_pack[590:586]);
    in_wt_norm[35] = cfg_is_fp16_d1[35] & (|in_wt_data_pack[574:570]);
    in_wt_norm[34] = cfg_is_fp16_d1[34] & (|in_wt_data_pack[558:554]);
    in_wt_norm[33] = cfg_is_fp16_d1[33] & (|in_wt_data_pack[542:538]);
    in_wt_norm[32] = cfg_is_fp16_d1[32] & (|in_wt_data_pack[526:522]);
    in_wt_norm[31] = cfg_is_fp16_d1[31] & (|in_wt_data_pack[510:506]);
    in_wt_norm[30] = cfg_is_fp16_d1[30] & (|in_wt_data_pack[494:490]);
    in_wt_norm[29] = cfg_is_fp16_d1[29] & (|in_wt_data_pack[478:474]);
    in_wt_norm[28] = cfg_is_fp16_d1[28] & (|in_wt_data_pack[462:458]);
    in_wt_norm[27] = cfg_is_fp16_d1[27] & (|in_wt_data_pack[446:442]);
    in_wt_norm[26] = cfg_is_fp16_d1[26] & (|in_wt_data_pack[430:426]);
    in_wt_norm[25] = cfg_is_fp16_d1[25] & (|in_wt_data_pack[414:410]);
    in_wt_norm[24] = cfg_is_fp16_d1[24] & (|in_wt_data_pack[398:394]);
    in_wt_norm[23] = cfg_is_fp16_d1[23] & (|in_wt_data_pack[382:378]);
    in_wt_norm[22] = cfg_is_fp16_d1[22] & (|in_wt_data_pack[366:362]);
    in_wt_norm[21] = cfg_is_fp16_d1[21] & (|in_wt_data_pack[350:346]);
    in_wt_norm[20] = cfg_is_fp16_d1[20] & (|in_wt_data_pack[334:330]);
    in_wt_norm[19] = cfg_is_fp16_d1[19] & (|in_wt_data_pack[318:314]);
    in_wt_norm[18] = cfg_is_fp16_d1[18] & (|in_wt_data_pack[302:298]);
    in_wt_norm[17] = cfg_is_fp16_d1[17] & (|in_wt_data_pack[286:282]);
    in_wt_norm[16] = cfg_is_fp16_d1[16] & (|in_wt_data_pack[270:266]);
    in_wt_norm[15] = cfg_is_fp16_d1[15] & (|in_wt_data_pack[254:250]);
    in_wt_norm[14] = cfg_is_fp16_d1[14] & (|in_wt_data_pack[238:234]);
    in_wt_norm[13] = cfg_is_fp16_d1[13] & (|in_wt_data_pack[222:218]);
    in_wt_norm[12] = cfg_is_fp16_d1[12] & (|in_wt_data_pack[206:202]);
    in_wt_norm[11] = cfg_is_fp16_d1[11] & (|in_wt_data_pack[190:186]);
    in_wt_norm[10] = cfg_is_fp16_d1[10] & (|in_wt_data_pack[174:170]);
    in_wt_norm[9] = cfg_is_fp16_d1[9] & (|in_wt_data_pack[158:154]);
    in_wt_norm[8] = cfg_is_fp16_d1[8] & (|in_wt_data_pack[142:138]);
    in_wt_norm[7] = cfg_is_fp16_d1[7] & (|in_wt_data_pack[126:122]);
    in_wt_norm[6] = cfg_is_fp16_d1[6] & (|in_wt_data_pack[110:106]);
    in_wt_norm[5] = cfg_is_fp16_d1[5] & (|in_wt_data_pack[94:90]);
    in_wt_norm[4] = cfg_is_fp16_d1[4] & (|in_wt_data_pack[78:74]);
    in_wt_norm[3] = cfg_is_fp16_d1[3] & (|in_wt_data_pack[62:58]);
    in_wt_norm[2] = cfg_is_fp16_d1[2] & (|in_wt_data_pack[46:42]);
    in_wt_norm[1] = cfg_is_fp16_d1[1] & (|in_wt_data_pack[30:26]);
    in_wt_norm[0] = cfg_is_fp16_d1[0] & (|in_wt_data_pack[14:10]);
end




always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori63 = ~cfg_is_fp16_d1[63] ? 12'b0 :
                                  in_wt_norm[63] ? {2'b1, in_wt_data_pack[1017:1008]} :
                                  {1'b0, in_wt_data_pack[1017:1008], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori62 = ~cfg_is_fp16_d1[62] ? 12'b0 :
                                  in_wt_norm[62] ? {2'b1, in_wt_data_pack[1001:992]} :
                                  {1'b0, in_wt_data_pack[1001:992], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori61 = ~cfg_is_fp16_d1[61] ? 12'b0 :
                                  in_wt_norm[61] ? {2'b1, in_wt_data_pack[985:976]} :
                                  {1'b0, in_wt_data_pack[985:976], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori60 = ~cfg_is_fp16_d1[60] ? 12'b0 :
                                  in_wt_norm[60] ? {2'b1, in_wt_data_pack[969:960]} :
                                  {1'b0, in_wt_data_pack[969:960], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori59 = ~cfg_is_fp16_d1[59] ? 12'b0 :
                                  in_wt_norm[59] ? {2'b1, in_wt_data_pack[953:944]} :
                                  {1'b0, in_wt_data_pack[953:944], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori58 = ~cfg_is_fp16_d1[58] ? 12'b0 :
                                  in_wt_norm[58] ? {2'b1, in_wt_data_pack[937:928]} :
                                  {1'b0, in_wt_data_pack[937:928], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori57 = ~cfg_is_fp16_d1[57] ? 12'b0 :
                                  in_wt_norm[57] ? {2'b1, in_wt_data_pack[921:912]} :
                                  {1'b0, in_wt_data_pack[921:912], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori56 = ~cfg_is_fp16_d1[56] ? 12'b0 :
                                  in_wt_norm[56] ? {2'b1, in_wt_data_pack[905:896]} :
                                  {1'b0, in_wt_data_pack[905:896], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori55 = ~cfg_is_fp16_d1[55] ? 12'b0 :
                                  in_wt_norm[55] ? {2'b1, in_wt_data_pack[889:880]} :
                                  {1'b0, in_wt_data_pack[889:880], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori54 = ~cfg_is_fp16_d1[54] ? 12'b0 :
                                  in_wt_norm[54] ? {2'b1, in_wt_data_pack[873:864]} :
                                  {1'b0, in_wt_data_pack[873:864], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori53 = ~cfg_is_fp16_d1[53] ? 12'b0 :
                                  in_wt_norm[53] ? {2'b1, in_wt_data_pack[857:848]} :
                                  {1'b0, in_wt_data_pack[857:848], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori52 = ~cfg_is_fp16_d1[52] ? 12'b0 :
                                  in_wt_norm[52] ? {2'b1, in_wt_data_pack[841:832]} :
                                  {1'b0, in_wt_data_pack[841:832], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori51 = ~cfg_is_fp16_d1[51] ? 12'b0 :
                                  in_wt_norm[51] ? {2'b1, in_wt_data_pack[825:816]} :
                                  {1'b0, in_wt_data_pack[825:816], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori50 = ~cfg_is_fp16_d1[50] ? 12'b0 :
                                  in_wt_norm[50] ? {2'b1, in_wt_data_pack[809:800]} :
                                  {1'b0, in_wt_data_pack[809:800], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori49 = ~cfg_is_fp16_d1[49] ? 12'b0 :
                                  in_wt_norm[49] ? {2'b1, in_wt_data_pack[793:784]} :
                                  {1'b0, in_wt_data_pack[793:784], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori48 = ~cfg_is_fp16_d1[48] ? 12'b0 :
                                  in_wt_norm[48] ? {2'b1, in_wt_data_pack[777:768]} :
                                  {1'b0, in_wt_data_pack[777:768], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori47 = ~cfg_is_fp16_d1[47] ? 12'b0 :
                                  in_wt_norm[47] ? {2'b1, in_wt_data_pack[761:752]} :
                                  {1'b0, in_wt_data_pack[761:752], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori46 = ~cfg_is_fp16_d1[46] ? 12'b0 :
                                  in_wt_norm[46] ? {2'b1, in_wt_data_pack[745:736]} :
                                  {1'b0, in_wt_data_pack[745:736], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori45 = ~cfg_is_fp16_d1[45] ? 12'b0 :
                                  in_wt_norm[45] ? {2'b1, in_wt_data_pack[729:720]} :
                                  {1'b0, in_wt_data_pack[729:720], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori44 = ~cfg_is_fp16_d1[44] ? 12'b0 :
                                  in_wt_norm[44] ? {2'b1, in_wt_data_pack[713:704]} :
                                  {1'b0, in_wt_data_pack[713:704], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori43 = ~cfg_is_fp16_d1[43] ? 12'b0 :
                                  in_wt_norm[43] ? {2'b1, in_wt_data_pack[697:688]} :
                                  {1'b0, in_wt_data_pack[697:688], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori42 = ~cfg_is_fp16_d1[42] ? 12'b0 :
                                  in_wt_norm[42] ? {2'b1, in_wt_data_pack[681:672]} :
                                  {1'b0, in_wt_data_pack[681:672], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori41 = ~cfg_is_fp16_d1[41] ? 12'b0 :
                                  in_wt_norm[41] ? {2'b1, in_wt_data_pack[665:656]} :
                                  {1'b0, in_wt_data_pack[665:656], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori40 = ~cfg_is_fp16_d1[40] ? 12'b0 :
                                  in_wt_norm[40] ? {2'b1, in_wt_data_pack[649:640]} :
                                  {1'b0, in_wt_data_pack[649:640], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori39 = ~cfg_is_fp16_d1[39] ? 12'b0 :
                                  in_wt_norm[39] ? {2'b1, in_wt_data_pack[633:624]} :
                                  {1'b0, in_wt_data_pack[633:624], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori38 = ~cfg_is_fp16_d1[38] ? 12'b0 :
                                  in_wt_norm[38] ? {2'b1, in_wt_data_pack[617:608]} :
                                  {1'b0, in_wt_data_pack[617:608], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori37 = ~cfg_is_fp16_d1[37] ? 12'b0 :
                                  in_wt_norm[37] ? {2'b1, in_wt_data_pack[601:592]} :
                                  {1'b0, in_wt_data_pack[601:592], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori36 = ~cfg_is_fp16_d1[36] ? 12'b0 :
                                  in_wt_norm[36] ? {2'b1, in_wt_data_pack[585:576]} :
                                  {1'b0, in_wt_data_pack[585:576], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori35 = ~cfg_is_fp16_d1[35] ? 12'b0 :
                                  in_wt_norm[35] ? {2'b1, in_wt_data_pack[569:560]} :
                                  {1'b0, in_wt_data_pack[569:560], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori34 = ~cfg_is_fp16_d1[34] ? 12'b0 :
                                  in_wt_norm[34] ? {2'b1, in_wt_data_pack[553:544]} :
                                  {1'b0, in_wt_data_pack[553:544], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori33 = ~cfg_is_fp16_d1[33] ? 12'b0 :
                                  in_wt_norm[33] ? {2'b1, in_wt_data_pack[537:528]} :
                                  {1'b0, in_wt_data_pack[537:528], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori32 = ~cfg_is_fp16_d1[32] ? 12'b0 :
                                  in_wt_norm[32] ? {2'b1, in_wt_data_pack[521:512]} :
                                  {1'b0, in_wt_data_pack[521:512], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori31 = ~cfg_is_fp16_d1[31] ? 12'b0 :
                                  in_wt_norm[31] ? {2'b1, in_wt_data_pack[505:496]} :
                                  {1'b0, in_wt_data_pack[505:496], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori30 = ~cfg_is_fp16_d1[30] ? 12'b0 :
                                  in_wt_norm[30] ? {2'b1, in_wt_data_pack[489:480]} :
                                  {1'b0, in_wt_data_pack[489:480], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori29 = ~cfg_is_fp16_d1[29] ? 12'b0 :
                                  in_wt_norm[29] ? {2'b1, in_wt_data_pack[473:464]} :
                                  {1'b0, in_wt_data_pack[473:464], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori28 = ~cfg_is_fp16_d1[28] ? 12'b0 :
                                  in_wt_norm[28] ? {2'b1, in_wt_data_pack[457:448]} :
                                  {1'b0, in_wt_data_pack[457:448], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori27 = ~cfg_is_fp16_d1[27] ? 12'b0 :
                                  in_wt_norm[27] ? {2'b1, in_wt_data_pack[441:432]} :
                                  {1'b0, in_wt_data_pack[441:432], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori26 = ~cfg_is_fp16_d1[26] ? 12'b0 :
                                  in_wt_norm[26] ? {2'b1, in_wt_data_pack[425:416]} :
                                  {1'b0, in_wt_data_pack[425:416], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori25 = ~cfg_is_fp16_d1[25] ? 12'b0 :
                                  in_wt_norm[25] ? {2'b1, in_wt_data_pack[409:400]} :
                                  {1'b0, in_wt_data_pack[409:400], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori24 = ~cfg_is_fp16_d1[24] ? 12'b0 :
                                  in_wt_norm[24] ? {2'b1, in_wt_data_pack[393:384]} :
                                  {1'b0, in_wt_data_pack[393:384], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori23 = ~cfg_is_fp16_d1[23] ? 12'b0 :
                                  in_wt_norm[23] ? {2'b1, in_wt_data_pack[377:368]} :
                                  {1'b0, in_wt_data_pack[377:368], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori22 = ~cfg_is_fp16_d1[22] ? 12'b0 :
                                  in_wt_norm[22] ? {2'b1, in_wt_data_pack[361:352]} :
                                  {1'b0, in_wt_data_pack[361:352], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori21 = ~cfg_is_fp16_d1[21] ? 12'b0 :
                                  in_wt_norm[21] ? {2'b1, in_wt_data_pack[345:336]} :
                                  {1'b0, in_wt_data_pack[345:336], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori20 = ~cfg_is_fp16_d1[20] ? 12'b0 :
                                  in_wt_norm[20] ? {2'b1, in_wt_data_pack[329:320]} :
                                  {1'b0, in_wt_data_pack[329:320], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori19 = ~cfg_is_fp16_d1[19] ? 12'b0 :
                                  in_wt_norm[19] ? {2'b1, in_wt_data_pack[313:304]} :
                                  {1'b0, in_wt_data_pack[313:304], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori18 = ~cfg_is_fp16_d1[18] ? 12'b0 :
                                  in_wt_norm[18] ? {2'b1, in_wt_data_pack[297:288]} :
                                  {1'b0, in_wt_data_pack[297:288], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori17 = ~cfg_is_fp16_d1[17] ? 12'b0 :
                                  in_wt_norm[17] ? {2'b1, in_wt_data_pack[281:272]} :
                                  {1'b0, in_wt_data_pack[281:272], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori16 = ~cfg_is_fp16_d1[16] ? 12'b0 :
                                  in_wt_norm[16] ? {2'b1, in_wt_data_pack[265:256]} :
                                  {1'b0, in_wt_data_pack[265:256], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori15 = ~cfg_is_fp16_d1[15] ? 12'b0 :
                                  in_wt_norm[15] ? {2'b1, in_wt_data_pack[249:240]} :
                                  {1'b0, in_wt_data_pack[249:240], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori14 = ~cfg_is_fp16_d1[14] ? 12'b0 :
                                  in_wt_norm[14] ? {2'b1, in_wt_data_pack[233:224]} :
                                  {1'b0, in_wt_data_pack[233:224], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori13 = ~cfg_is_fp16_d1[13] ? 12'b0 :
                                  in_wt_norm[13] ? {2'b1, in_wt_data_pack[217:208]} :
                                  {1'b0, in_wt_data_pack[217:208], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori12 = ~cfg_is_fp16_d1[12] ? 12'b0 :
                                  in_wt_norm[12] ? {2'b1, in_wt_data_pack[201:192]} :
                                  {1'b0, in_wt_data_pack[201:192], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori11 = ~cfg_is_fp16_d1[11] ? 12'b0 :
                                  in_wt_norm[11] ? {2'b1, in_wt_data_pack[185:176]} :
                                  {1'b0, in_wt_data_pack[185:176], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori10 = ~cfg_is_fp16_d1[10] ? 12'b0 :
                                  in_wt_norm[10] ? {2'b1, in_wt_data_pack[169:160]} :
                                  {1'b0, in_wt_data_pack[169:160], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori9 = ~cfg_is_fp16_d1[9] ? 12'b0 :
                                  in_wt_norm[9] ? {2'b1, in_wt_data_pack[153:144]} :
                                  {1'b0, in_wt_data_pack[153:144], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori8 = ~cfg_is_fp16_d1[8] ? 12'b0 :
                                  in_wt_norm[8] ? {2'b1, in_wt_data_pack[137:128]} :
                                  {1'b0, in_wt_data_pack[137:128], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori7 = ~cfg_is_fp16_d1[7] ? 12'b0 :
                                  in_wt_norm[7] ? {2'b1, in_wt_data_pack[121:112]} :
                                  {1'b0, in_wt_data_pack[121:112], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori6 = ~cfg_is_fp16_d1[6] ? 12'b0 :
                                  in_wt_norm[6] ? {2'b1, in_wt_data_pack[105:96]} :
                                  {1'b0, in_wt_data_pack[105:96], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori5 = ~cfg_is_fp16_d1[5] ? 12'b0 :
                                  in_wt_norm[5] ? {2'b1, in_wt_data_pack[89:80]} :
                                  {1'b0, in_wt_data_pack[89:80], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori4 = ~cfg_is_fp16_d1[4] ? 12'b0 :
                                  in_wt_norm[4] ? {2'b1, in_wt_data_pack[73:64]} :
                                  {1'b0, in_wt_data_pack[73:64], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori3 = ~cfg_is_fp16_d1[3] ? 12'b0 :
                                  in_wt_norm[3] ? {2'b1, in_wt_data_pack[57:48]} :
                                  {1'b0, in_wt_data_pack[57:48], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori2 = ~cfg_is_fp16_d1[2] ? 12'b0 :
                                  in_wt_norm[2] ? {2'b1, in_wt_data_pack[41:32]} :
                                  {1'b0, in_wt_data_pack[41:32], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori1 = ~cfg_is_fp16_d1[1] ? 12'b0 :
                                  in_wt_norm[1] ? {2'b1, in_wt_data_pack[25:16]} :
                                  {1'b0, in_wt_data_pack[25:16], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_wt_norm
  or in_wt_data_pack
  ) begin
    in_wt_data_fp16_mts_ori0 = ~cfg_is_fp16_d1[0] ? 12'b0 :
                                  in_wt_norm[0] ? {2'b1, in_wt_data_pack[9:0]} :
                                  {1'b0, in_wt_data_pack[9:0], 1'b0};
end







always @(
  in_wt_data_fp16_mts_ori63
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft63[14:0] = ({3'b0, in_wt_data_fp16_mts_ori63} << in_wt_data_pack[1019:1018]);
    in_wt_data_fp16_63 = ({16{cfg_is_fp16_d1[63]}} & {in_wt_data_pack[1023], in_wt_data_fp16_mts_sft63});
end



always @(
  in_wt_data_fp16_mts_ori62
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft62[14:0] = ({3'b0, in_wt_data_fp16_mts_ori62} << in_wt_data_pack[1003:1002]);
    in_wt_data_fp16_62 = ({16{cfg_is_fp16_d1[62]}} & {in_wt_data_pack[1007], in_wt_data_fp16_mts_sft62});
end



always @(
  in_wt_data_fp16_mts_ori61
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft61[14:0] = ({3'b0, in_wt_data_fp16_mts_ori61} << in_wt_data_pack[987:986]);
    in_wt_data_fp16_61 = ({16{cfg_is_fp16_d1[61]}} & {in_wt_data_pack[991], in_wt_data_fp16_mts_sft61});
end



always @(
  in_wt_data_fp16_mts_ori60
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft60[14:0] = ({3'b0, in_wt_data_fp16_mts_ori60} << in_wt_data_pack[971:970]);
    in_wt_data_fp16_60 = ({16{cfg_is_fp16_d1[60]}} & {in_wt_data_pack[975], in_wt_data_fp16_mts_sft60});
end



always @(
  in_wt_data_fp16_mts_ori59
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft59[14:0] = ({3'b0, in_wt_data_fp16_mts_ori59} << in_wt_data_pack[955:954]);
    in_wt_data_fp16_59 = ({16{cfg_is_fp16_d1[59]}} & {in_wt_data_pack[959], in_wt_data_fp16_mts_sft59});
end



always @(
  in_wt_data_fp16_mts_ori58
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft58[14:0] = ({3'b0, in_wt_data_fp16_mts_ori58} << in_wt_data_pack[939:938]);
    in_wt_data_fp16_58 = ({16{cfg_is_fp16_d1[58]}} & {in_wt_data_pack[943], in_wt_data_fp16_mts_sft58});
end



always @(
  in_wt_data_fp16_mts_ori57
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft57[14:0] = ({3'b0, in_wt_data_fp16_mts_ori57} << in_wt_data_pack[923:922]);
    in_wt_data_fp16_57 = ({16{cfg_is_fp16_d1[57]}} & {in_wt_data_pack[927], in_wt_data_fp16_mts_sft57});
end



always @(
  in_wt_data_fp16_mts_ori56
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft56[14:0] = ({3'b0, in_wt_data_fp16_mts_ori56} << in_wt_data_pack[907:906]);
    in_wt_data_fp16_56 = ({16{cfg_is_fp16_d1[56]}} & {in_wt_data_pack[911], in_wt_data_fp16_mts_sft56});
end



always @(
  in_wt_data_fp16_mts_ori55
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft55[14:0] = ({3'b0, in_wt_data_fp16_mts_ori55} << in_wt_data_pack[891:890]);
    in_wt_data_fp16_55 = ({16{cfg_is_fp16_d1[55]}} & {in_wt_data_pack[895], in_wt_data_fp16_mts_sft55});
end



always @(
  in_wt_data_fp16_mts_ori54
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft54[14:0] = ({3'b0, in_wt_data_fp16_mts_ori54} << in_wt_data_pack[875:874]);
    in_wt_data_fp16_54 = ({16{cfg_is_fp16_d1[54]}} & {in_wt_data_pack[879], in_wt_data_fp16_mts_sft54});
end



always @(
  in_wt_data_fp16_mts_ori53
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft53[14:0] = ({3'b0, in_wt_data_fp16_mts_ori53} << in_wt_data_pack[859:858]);
    in_wt_data_fp16_53 = ({16{cfg_is_fp16_d1[53]}} & {in_wt_data_pack[863], in_wt_data_fp16_mts_sft53});
end



always @(
  in_wt_data_fp16_mts_ori52
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft52[14:0] = ({3'b0, in_wt_data_fp16_mts_ori52} << in_wt_data_pack[843:842]);
    in_wt_data_fp16_52 = ({16{cfg_is_fp16_d1[52]}} & {in_wt_data_pack[847], in_wt_data_fp16_mts_sft52});
end



always @(
  in_wt_data_fp16_mts_ori51
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft51[14:0] = ({3'b0, in_wt_data_fp16_mts_ori51} << in_wt_data_pack[827:826]);
    in_wt_data_fp16_51 = ({16{cfg_is_fp16_d1[51]}} & {in_wt_data_pack[831], in_wt_data_fp16_mts_sft51});
end



always @(
  in_wt_data_fp16_mts_ori50
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft50[14:0] = ({3'b0, in_wt_data_fp16_mts_ori50} << in_wt_data_pack[811:810]);
    in_wt_data_fp16_50 = ({16{cfg_is_fp16_d1[50]}} & {in_wt_data_pack[815], in_wt_data_fp16_mts_sft50});
end



always @(
  in_wt_data_fp16_mts_ori49
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft49[14:0] = ({3'b0, in_wt_data_fp16_mts_ori49} << in_wt_data_pack[795:794]);
    in_wt_data_fp16_49 = ({16{cfg_is_fp16_d1[49]}} & {in_wt_data_pack[799], in_wt_data_fp16_mts_sft49});
end



always @(
  in_wt_data_fp16_mts_ori48
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft48[14:0] = ({3'b0, in_wt_data_fp16_mts_ori48} << in_wt_data_pack[779:778]);
    in_wt_data_fp16_48 = ({16{cfg_is_fp16_d1[48]}} & {in_wt_data_pack[783], in_wt_data_fp16_mts_sft48});
end



always @(
  in_wt_data_fp16_mts_ori47
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft47[14:0] = ({3'b0, in_wt_data_fp16_mts_ori47} << in_wt_data_pack[763:762]);
    in_wt_data_fp16_47 = ({16{cfg_is_fp16_d1[47]}} & {in_wt_data_pack[767], in_wt_data_fp16_mts_sft47});
end



always @(
  in_wt_data_fp16_mts_ori46
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft46[14:0] = ({3'b0, in_wt_data_fp16_mts_ori46} << in_wt_data_pack[747:746]);
    in_wt_data_fp16_46 = ({16{cfg_is_fp16_d1[46]}} & {in_wt_data_pack[751], in_wt_data_fp16_mts_sft46});
end



always @(
  in_wt_data_fp16_mts_ori45
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft45[14:0] = ({3'b0, in_wt_data_fp16_mts_ori45} << in_wt_data_pack[731:730]);
    in_wt_data_fp16_45 = ({16{cfg_is_fp16_d1[45]}} & {in_wt_data_pack[735], in_wt_data_fp16_mts_sft45});
end



always @(
  in_wt_data_fp16_mts_ori44
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft44[14:0] = ({3'b0, in_wt_data_fp16_mts_ori44} << in_wt_data_pack[715:714]);
    in_wt_data_fp16_44 = ({16{cfg_is_fp16_d1[44]}} & {in_wt_data_pack[719], in_wt_data_fp16_mts_sft44});
end



always @(
  in_wt_data_fp16_mts_ori43
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft43[14:0] = ({3'b0, in_wt_data_fp16_mts_ori43} << in_wt_data_pack[699:698]);
    in_wt_data_fp16_43 = ({16{cfg_is_fp16_d1[43]}} & {in_wt_data_pack[703], in_wt_data_fp16_mts_sft43});
end



always @(
  in_wt_data_fp16_mts_ori42
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft42[14:0] = ({3'b0, in_wt_data_fp16_mts_ori42} << in_wt_data_pack[683:682]);
    in_wt_data_fp16_42 = ({16{cfg_is_fp16_d1[42]}} & {in_wt_data_pack[687], in_wt_data_fp16_mts_sft42});
end



always @(
  in_wt_data_fp16_mts_ori41
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft41[14:0] = ({3'b0, in_wt_data_fp16_mts_ori41} << in_wt_data_pack[667:666]);
    in_wt_data_fp16_41 = ({16{cfg_is_fp16_d1[41]}} & {in_wt_data_pack[671], in_wt_data_fp16_mts_sft41});
end



always @(
  in_wt_data_fp16_mts_ori40
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft40[14:0] = ({3'b0, in_wt_data_fp16_mts_ori40} << in_wt_data_pack[651:650]);
    in_wt_data_fp16_40 = ({16{cfg_is_fp16_d1[40]}} & {in_wt_data_pack[655], in_wt_data_fp16_mts_sft40});
end



always @(
  in_wt_data_fp16_mts_ori39
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft39[14:0] = ({3'b0, in_wt_data_fp16_mts_ori39} << in_wt_data_pack[635:634]);
    in_wt_data_fp16_39 = ({16{cfg_is_fp16_d1[39]}} & {in_wt_data_pack[639], in_wt_data_fp16_mts_sft39});
end



always @(
  in_wt_data_fp16_mts_ori38
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft38[14:0] = ({3'b0, in_wt_data_fp16_mts_ori38} << in_wt_data_pack[619:618]);
    in_wt_data_fp16_38 = ({16{cfg_is_fp16_d1[38]}} & {in_wt_data_pack[623], in_wt_data_fp16_mts_sft38});
end



always @(
  in_wt_data_fp16_mts_ori37
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft37[14:0] = ({3'b0, in_wt_data_fp16_mts_ori37} << in_wt_data_pack[603:602]);
    in_wt_data_fp16_37 = ({16{cfg_is_fp16_d1[37]}} & {in_wt_data_pack[607], in_wt_data_fp16_mts_sft37});
end



always @(
  in_wt_data_fp16_mts_ori36
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft36[14:0] = ({3'b0, in_wt_data_fp16_mts_ori36} << in_wt_data_pack[587:586]);
    in_wt_data_fp16_36 = ({16{cfg_is_fp16_d1[36]}} & {in_wt_data_pack[591], in_wt_data_fp16_mts_sft36});
end



always @(
  in_wt_data_fp16_mts_ori35
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft35[14:0] = ({3'b0, in_wt_data_fp16_mts_ori35} << in_wt_data_pack[571:570]);
    in_wt_data_fp16_35 = ({16{cfg_is_fp16_d1[35]}} & {in_wt_data_pack[575], in_wt_data_fp16_mts_sft35});
end



always @(
  in_wt_data_fp16_mts_ori34
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft34[14:0] = ({3'b0, in_wt_data_fp16_mts_ori34} << in_wt_data_pack[555:554]);
    in_wt_data_fp16_34 = ({16{cfg_is_fp16_d1[34]}} & {in_wt_data_pack[559], in_wt_data_fp16_mts_sft34});
end



always @(
  in_wt_data_fp16_mts_ori33
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft33[14:0] = ({3'b0, in_wt_data_fp16_mts_ori33} << in_wt_data_pack[539:538]);
    in_wt_data_fp16_33 = ({16{cfg_is_fp16_d1[33]}} & {in_wt_data_pack[543], in_wt_data_fp16_mts_sft33});
end



always @(
  in_wt_data_fp16_mts_ori32
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft32[14:0] = ({3'b0, in_wt_data_fp16_mts_ori32} << in_wt_data_pack[523:522]);
    in_wt_data_fp16_32 = ({16{cfg_is_fp16_d1[32]}} & {in_wt_data_pack[527], in_wt_data_fp16_mts_sft32});
end



always @(
  in_wt_data_fp16_mts_ori31
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft31[14:0] = ({3'b0, in_wt_data_fp16_mts_ori31} << in_wt_data_pack[507:506]);
    in_wt_data_fp16_31 = ({16{cfg_is_fp16_d1[31]}} & {in_wt_data_pack[511], in_wt_data_fp16_mts_sft31});
end



always @(
  in_wt_data_fp16_mts_ori30
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft30[14:0] = ({3'b0, in_wt_data_fp16_mts_ori30} << in_wt_data_pack[491:490]);
    in_wt_data_fp16_30 = ({16{cfg_is_fp16_d1[30]}} & {in_wt_data_pack[495], in_wt_data_fp16_mts_sft30});
end



always @(
  in_wt_data_fp16_mts_ori29
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft29[14:0] = ({3'b0, in_wt_data_fp16_mts_ori29} << in_wt_data_pack[475:474]);
    in_wt_data_fp16_29 = ({16{cfg_is_fp16_d1[29]}} & {in_wt_data_pack[479], in_wt_data_fp16_mts_sft29});
end



always @(
  in_wt_data_fp16_mts_ori28
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft28[14:0] = ({3'b0, in_wt_data_fp16_mts_ori28} << in_wt_data_pack[459:458]);
    in_wt_data_fp16_28 = ({16{cfg_is_fp16_d1[28]}} & {in_wt_data_pack[463], in_wt_data_fp16_mts_sft28});
end



always @(
  in_wt_data_fp16_mts_ori27
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft27[14:0] = ({3'b0, in_wt_data_fp16_mts_ori27} << in_wt_data_pack[443:442]);
    in_wt_data_fp16_27 = ({16{cfg_is_fp16_d1[27]}} & {in_wt_data_pack[447], in_wt_data_fp16_mts_sft27});
end



always @(
  in_wt_data_fp16_mts_ori26
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft26[14:0] = ({3'b0, in_wt_data_fp16_mts_ori26} << in_wt_data_pack[427:426]);
    in_wt_data_fp16_26 = ({16{cfg_is_fp16_d1[26]}} & {in_wt_data_pack[431], in_wt_data_fp16_mts_sft26});
end



always @(
  in_wt_data_fp16_mts_ori25
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft25[14:0] = ({3'b0, in_wt_data_fp16_mts_ori25} << in_wt_data_pack[411:410]);
    in_wt_data_fp16_25 = ({16{cfg_is_fp16_d1[25]}} & {in_wt_data_pack[415], in_wt_data_fp16_mts_sft25});
end



always @(
  in_wt_data_fp16_mts_ori24
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft24[14:0] = ({3'b0, in_wt_data_fp16_mts_ori24} << in_wt_data_pack[395:394]);
    in_wt_data_fp16_24 = ({16{cfg_is_fp16_d1[24]}} & {in_wt_data_pack[399], in_wt_data_fp16_mts_sft24});
end



always @(
  in_wt_data_fp16_mts_ori23
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft23[14:0] = ({3'b0, in_wt_data_fp16_mts_ori23} << in_wt_data_pack[379:378]);
    in_wt_data_fp16_23 = ({16{cfg_is_fp16_d1[23]}} & {in_wt_data_pack[383], in_wt_data_fp16_mts_sft23});
end



always @(
  in_wt_data_fp16_mts_ori22
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft22[14:0] = ({3'b0, in_wt_data_fp16_mts_ori22} << in_wt_data_pack[363:362]);
    in_wt_data_fp16_22 = ({16{cfg_is_fp16_d1[22]}} & {in_wt_data_pack[367], in_wt_data_fp16_mts_sft22});
end



always @(
  in_wt_data_fp16_mts_ori21
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft21[14:0] = ({3'b0, in_wt_data_fp16_mts_ori21} << in_wt_data_pack[347:346]);
    in_wt_data_fp16_21 = ({16{cfg_is_fp16_d1[21]}} & {in_wt_data_pack[351], in_wt_data_fp16_mts_sft21});
end



always @(
  in_wt_data_fp16_mts_ori20
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft20[14:0] = ({3'b0, in_wt_data_fp16_mts_ori20} << in_wt_data_pack[331:330]);
    in_wt_data_fp16_20 = ({16{cfg_is_fp16_d1[20]}} & {in_wt_data_pack[335], in_wt_data_fp16_mts_sft20});
end



always @(
  in_wt_data_fp16_mts_ori19
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft19[14:0] = ({3'b0, in_wt_data_fp16_mts_ori19} << in_wt_data_pack[315:314]);
    in_wt_data_fp16_19 = ({16{cfg_is_fp16_d1[19]}} & {in_wt_data_pack[319], in_wt_data_fp16_mts_sft19});
end



always @(
  in_wt_data_fp16_mts_ori18
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft18[14:0] = ({3'b0, in_wt_data_fp16_mts_ori18} << in_wt_data_pack[299:298]);
    in_wt_data_fp16_18 = ({16{cfg_is_fp16_d1[18]}} & {in_wt_data_pack[303], in_wt_data_fp16_mts_sft18});
end



always @(
  in_wt_data_fp16_mts_ori17
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft17[14:0] = ({3'b0, in_wt_data_fp16_mts_ori17} << in_wt_data_pack[283:282]);
    in_wt_data_fp16_17 = ({16{cfg_is_fp16_d1[17]}} & {in_wt_data_pack[287], in_wt_data_fp16_mts_sft17});
end



always @(
  in_wt_data_fp16_mts_ori16
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft16[14:0] = ({3'b0, in_wt_data_fp16_mts_ori16} << in_wt_data_pack[267:266]);
    in_wt_data_fp16_16 = ({16{cfg_is_fp16_d1[16]}} & {in_wt_data_pack[271], in_wt_data_fp16_mts_sft16});
end



always @(
  in_wt_data_fp16_mts_ori15
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft15[14:0] = ({3'b0, in_wt_data_fp16_mts_ori15} << in_wt_data_pack[251:250]);
    in_wt_data_fp16_15 = ({16{cfg_is_fp16_d1[15]}} & {in_wt_data_pack[255], in_wt_data_fp16_mts_sft15});
end



always @(
  in_wt_data_fp16_mts_ori14
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft14[14:0] = ({3'b0, in_wt_data_fp16_mts_ori14} << in_wt_data_pack[235:234]);
    in_wt_data_fp16_14 = ({16{cfg_is_fp16_d1[14]}} & {in_wt_data_pack[239], in_wt_data_fp16_mts_sft14});
end



always @(
  in_wt_data_fp16_mts_ori13
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft13[14:0] = ({3'b0, in_wt_data_fp16_mts_ori13} << in_wt_data_pack[219:218]);
    in_wt_data_fp16_13 = ({16{cfg_is_fp16_d1[13]}} & {in_wt_data_pack[223], in_wt_data_fp16_mts_sft13});
end



always @(
  in_wt_data_fp16_mts_ori12
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft12[14:0] = ({3'b0, in_wt_data_fp16_mts_ori12} << in_wt_data_pack[203:202]);
    in_wt_data_fp16_12 = ({16{cfg_is_fp16_d1[12]}} & {in_wt_data_pack[207], in_wt_data_fp16_mts_sft12});
end



always @(
  in_wt_data_fp16_mts_ori11
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft11[14:0] = ({3'b0, in_wt_data_fp16_mts_ori11} << in_wt_data_pack[187:186]);
    in_wt_data_fp16_11 = ({16{cfg_is_fp16_d1[11]}} & {in_wt_data_pack[191], in_wt_data_fp16_mts_sft11});
end



always @(
  in_wt_data_fp16_mts_ori10
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft10[14:0] = ({3'b0, in_wt_data_fp16_mts_ori10} << in_wt_data_pack[171:170]);
    in_wt_data_fp16_10 = ({16{cfg_is_fp16_d1[10]}} & {in_wt_data_pack[175], in_wt_data_fp16_mts_sft10});
end



always @(
  in_wt_data_fp16_mts_ori9
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft9[14:0] = ({3'b0, in_wt_data_fp16_mts_ori9} << in_wt_data_pack[155:154]);
    in_wt_data_fp16_9 = ({16{cfg_is_fp16_d1[9]}} & {in_wt_data_pack[159], in_wt_data_fp16_mts_sft9});
end



always @(
  in_wt_data_fp16_mts_ori8
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft8[14:0] = ({3'b0, in_wt_data_fp16_mts_ori8} << in_wt_data_pack[139:138]);
    in_wt_data_fp16_8 = ({16{cfg_is_fp16_d1[8]}} & {in_wt_data_pack[143], in_wt_data_fp16_mts_sft8});
end



always @(
  in_wt_data_fp16_mts_ori7
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft7[14:0] = ({3'b0, in_wt_data_fp16_mts_ori7} << in_wt_data_pack[123:122]);
    in_wt_data_fp16_7 = ({16{cfg_is_fp16_d1[7]}} & {in_wt_data_pack[127], in_wt_data_fp16_mts_sft7});
end



always @(
  in_wt_data_fp16_mts_ori6
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft6[14:0] = ({3'b0, in_wt_data_fp16_mts_ori6} << in_wt_data_pack[107:106]);
    in_wt_data_fp16_6 = ({16{cfg_is_fp16_d1[6]}} & {in_wt_data_pack[111], in_wt_data_fp16_mts_sft6});
end



always @(
  in_wt_data_fp16_mts_ori5
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft5[14:0] = ({3'b0, in_wt_data_fp16_mts_ori5} << in_wt_data_pack[91:90]);
    in_wt_data_fp16_5 = ({16{cfg_is_fp16_d1[5]}} & {in_wt_data_pack[95], in_wt_data_fp16_mts_sft5});
end



always @(
  in_wt_data_fp16_mts_ori4
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft4[14:0] = ({3'b0, in_wt_data_fp16_mts_ori4} << in_wt_data_pack[75:74]);
    in_wt_data_fp16_4 = ({16{cfg_is_fp16_d1[4]}} & {in_wt_data_pack[79], in_wt_data_fp16_mts_sft4});
end



always @(
  in_wt_data_fp16_mts_ori3
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft3[14:0] = ({3'b0, in_wt_data_fp16_mts_ori3} << in_wt_data_pack[59:58]);
    in_wt_data_fp16_3 = ({16{cfg_is_fp16_d1[3]}} & {in_wt_data_pack[63], in_wt_data_fp16_mts_sft3});
end



always @(
  in_wt_data_fp16_mts_ori2
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft2[14:0] = ({3'b0, in_wt_data_fp16_mts_ori2} << in_wt_data_pack[43:42]);
    in_wt_data_fp16_2 = ({16{cfg_is_fp16_d1[2]}} & {in_wt_data_pack[47], in_wt_data_fp16_mts_sft2});
end



always @(
  in_wt_data_fp16_mts_ori1
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft1[14:0] = ({3'b0, in_wt_data_fp16_mts_ori1} << in_wt_data_pack[27:26]);
    in_wt_data_fp16_1 = ({16{cfg_is_fp16_d1[1]}} & {in_wt_data_pack[31], in_wt_data_fp16_mts_sft1});
end



always @(
  in_wt_data_fp16_mts_ori0
  or in_wt_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_wt_data_fp16_mts_sft0[14:0] = ({3'b0, in_wt_data_fp16_mts_ori0} << in_wt_data_pack[11:10]);
    in_wt_data_fp16_0 = ({16{cfg_is_fp16_d1[0]}} & {in_wt_data_pack[15], in_wt_data_fp16_mts_sft0});
end







always @(
  in_wt_nan
  ) begin
    wt_has_nan = (|in_wt_nan);
end

always @(
  in_wt_data_fp16_63
  or in_wt_data_fp16_62
  or in_wt_data_fp16_61
  or in_wt_data_fp16_60
  or in_wt_data_fp16_59
  or in_wt_data_fp16_58
  or in_wt_data_fp16_57
  or in_wt_data_fp16_56
  or in_wt_data_fp16_55
  or in_wt_data_fp16_54
  or in_wt_data_fp16_53
  or in_wt_data_fp16_52
  or in_wt_data_fp16_51
  or in_wt_data_fp16_50
  or in_wt_data_fp16_49
  or in_wt_data_fp16_48
  or in_wt_data_fp16_47
  or in_wt_data_fp16_46
  or in_wt_data_fp16_45
  or in_wt_data_fp16_44
  or in_wt_data_fp16_43
  or in_wt_data_fp16_42
  or in_wt_data_fp16_41
  or in_wt_data_fp16_40
  or in_wt_data_fp16_39
  or in_wt_data_fp16_38
  or in_wt_data_fp16_37
  or in_wt_data_fp16_36
  or in_wt_data_fp16_35
  or in_wt_data_fp16_34
  or in_wt_data_fp16_33
  or in_wt_data_fp16_32
  or in_wt_data_fp16_31
  or in_wt_data_fp16_30
  or in_wt_data_fp16_29
  or in_wt_data_fp16_28
  or in_wt_data_fp16_27
  or in_wt_data_fp16_26
  or in_wt_data_fp16_25
  or in_wt_data_fp16_24
  or in_wt_data_fp16_23
  or in_wt_data_fp16_22
  or in_wt_data_fp16_21
  or in_wt_data_fp16_20
  or in_wt_data_fp16_19
  or in_wt_data_fp16_18
  or in_wt_data_fp16_17
  or in_wt_data_fp16_16
  or in_wt_data_fp16_15
  or in_wt_data_fp16_14
  or in_wt_data_fp16_13
  or in_wt_data_fp16_12
  or in_wt_data_fp16_11
  or in_wt_data_fp16_10
  or in_wt_data_fp16_9
  or in_wt_data_fp16_8
  or in_wt_data_fp16_7
  or in_wt_data_fp16_6
  or in_wt_data_fp16_5
  or in_wt_data_fp16_4
  or in_wt_data_fp16_3
  or in_wt_data_fp16_2
  or in_wt_data_fp16_1
  or in_wt_data_fp16_0
  ) begin
    in_wt_data_fp16 = {in_wt_data_fp16_63, in_wt_data_fp16_62, in_wt_data_fp16_61, in_wt_data_fp16_60, in_wt_data_fp16_59, in_wt_data_fp16_58, in_wt_data_fp16_57, in_wt_data_fp16_56, in_wt_data_fp16_55, in_wt_data_fp16_54, in_wt_data_fp16_53, in_wt_data_fp16_52, in_wt_data_fp16_51, in_wt_data_fp16_50, in_wt_data_fp16_49, in_wt_data_fp16_48, in_wt_data_fp16_47, in_wt_data_fp16_46, in_wt_data_fp16_45, in_wt_data_fp16_44, in_wt_data_fp16_43, in_wt_data_fp16_42, in_wt_data_fp16_41, in_wt_data_fp16_40, in_wt_data_fp16_39, in_wt_data_fp16_38, in_wt_data_fp16_37, in_wt_data_fp16_36, in_wt_data_fp16_35, in_wt_data_fp16_34, in_wt_data_fp16_33, in_wt_data_fp16_32, in_wt_data_fp16_31, in_wt_data_fp16_30, in_wt_data_fp16_29, in_wt_data_fp16_28, in_wt_data_fp16_27, in_wt_data_fp16_26, in_wt_data_fp16_25, in_wt_data_fp16_24, in_wt_data_fp16_23, in_wt_data_fp16_22, in_wt_data_fp16_21, in_wt_data_fp16_20, in_wt_data_fp16_19, in_wt_data_fp16_18, in_wt_data_fp16_17, in_wt_data_fp16_16, in_wt_data_fp16_15, in_wt_data_fp16_14, in_wt_data_fp16_13, in_wt_data_fp16_12, in_wt_data_fp16_11, in_wt_data_fp16_10, in_wt_data_fp16_9, in_wt_data_fp16_8, in_wt_data_fp16_7, in_wt_data_fp16_6, in_wt_data_fp16_5, in_wt_data_fp16_4, in_wt_data_fp16_3, in_wt_data_fp16_2, in_wt_data_fp16_1, in_wt_data_fp16_0};
end

//////////////// wt_pre_data_w ////////////////
always @(
  in_wt_data_fp16
  or in_wt_data_int8
  or in_wt_data_int16
  ) begin
    wt_pre_data_w = in_wt_data_fp16 | in_wt_data_int8 | in_wt_data_int16;
end

always @(
  cfg_is_fp16_d1
  or wt_has_nan
  or in_wt_mask
  or cfg_is_int8_d1
  or in_wt_mask_int8
  ) begin
    wt_pre_nz_w = (cfg_is_fp16_d1[64]) ? {128{~wt_has_nan}} & in_wt_mask :
                  (cfg_is_int8_d1[64]) ? in_wt_mask_int8 :
                  in_wt_mask;
end

always @(
  in_wt_exp
  ) begin
    wt_pre_exp_w = in_wt_exp;
end

always @(
  wt_pre_nz_w
  ) begin
    wt_pre_mask_w = {wt_pre_nz_w[63*2],wt_pre_nz_w[62*2],wt_pre_nz_w[61*2],wt_pre_nz_w[60*2],wt_pre_nz_w[59*2],wt_pre_nz_w[58*2],wt_pre_nz_w[57*2],wt_pre_nz_w[56*2],wt_pre_nz_w[55*2],wt_pre_nz_w[54*2],wt_pre_nz_w[53*2],wt_pre_nz_w[52*2],wt_pre_nz_w[51*2],wt_pre_nz_w[50*2],wt_pre_nz_w[49*2],wt_pre_nz_w[48*2],wt_pre_nz_w[47*2],wt_pre_nz_w[46*2],wt_pre_nz_w[45*2],wt_pre_nz_w[44*2],wt_pre_nz_w[43*2],wt_pre_nz_w[42*2],wt_pre_nz_w[41*2],wt_pre_nz_w[40*2],wt_pre_nz_w[39*2],wt_pre_nz_w[38*2],wt_pre_nz_w[37*2],wt_pre_nz_w[36*2],wt_pre_nz_w[35*2],wt_pre_nz_w[34*2],wt_pre_nz_w[33*2],wt_pre_nz_w[32*2],wt_pre_nz_w[31*2],wt_pre_nz_w[30*2],wt_pre_nz_w[29*2],wt_pre_nz_w[28*2],wt_pre_nz_w[27*2],wt_pre_nz_w[26*2],wt_pre_nz_w[25*2],wt_pre_nz_w[24*2],wt_pre_nz_w[23*2],wt_pre_nz_w[22*2],wt_pre_nz_w[21*2],wt_pre_nz_w[20*2],wt_pre_nz_w[19*2],wt_pre_nz_w[18*2],wt_pre_nz_w[17*2],wt_pre_nz_w[16*2],wt_pre_nz_w[15*2],wt_pre_nz_w[14*2],wt_pre_nz_w[13*2],wt_pre_nz_w[12*2],wt_pre_nz_w[11*2],wt_pre_nz_w[10*2],wt_pre_nz_w[9*2],wt_pre_nz_w[8*2],wt_pre_nz_w[7*2],wt_pre_nz_w[6*2],wt_pre_nz_w[5*2],wt_pre_nz_w[4*2],wt_pre_nz_w[3*2],wt_pre_nz_w[2*2],wt_pre_nz_w[1*2],wt_pre_nz_w[0*2]};
end

//==========================================================
// Weight pre-process register         
//==========================================================
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt_pre_sel <= {8{1'b0}};
  end else begin
  wt_pre_sel <= in_wt_sel;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld) == 1'b1) begin
    wt_pre_nz <= wt_pre_nz_w;
  // VCS coverage off
  end else if ((in_wt_pvld) == 1'b0) begin
  end else begin
    wt_pre_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b1) begin
    wt_pre_mask <= wt_pre_mask_w;
  // VCS coverage off
  end else if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b0) begin
  end else begin
    wt_pre_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b1) begin
    wt_pre_exp <= wt_pre_exp_w;
  // VCS coverage off
  end else if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b0) begin
  end else begin
    wt_pre_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b1) begin
    wt_pre_nan <= in_wt_nan;
  // VCS coverage off
  end else if ((in_wt_pvld & cfg_is_fp16_d1[65]) == 1'b0) begin
  end else begin
    wt_pre_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[0] | in_wt_nan[0])) == 1'b1) begin
    wt_pre_data[7:0] <= wt_pre_data_w[7:0];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[0] | in_wt_nan[0])) == 1'b0) begin
  end else begin
    wt_pre_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[1] | in_wt_nan[0])) == 1'b1) begin
    wt_pre_data[15:8] <= wt_pre_data_w[15:8];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[1] | in_wt_nan[0])) == 1'b0) begin
  end else begin
    wt_pre_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[2] | in_wt_nan[1])) == 1'b1) begin
    wt_pre_data[23:16] <= wt_pre_data_w[23:16];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[2] | in_wt_nan[1])) == 1'b0) begin
  end else begin
    wt_pre_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[3] | in_wt_nan[1])) == 1'b1) begin
    wt_pre_data[31:24] <= wt_pre_data_w[31:24];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[3] | in_wt_nan[1])) == 1'b0) begin
  end else begin
    wt_pre_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[4] | in_wt_nan[2])) == 1'b1) begin
    wt_pre_data[39:32] <= wt_pre_data_w[39:32];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[4] | in_wt_nan[2])) == 1'b0) begin
  end else begin
    wt_pre_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[5] | in_wt_nan[2])) == 1'b1) begin
    wt_pre_data[47:40] <= wt_pre_data_w[47:40];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[5] | in_wt_nan[2])) == 1'b0) begin
  end else begin
    wt_pre_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[6] | in_wt_nan[3])) == 1'b1) begin
    wt_pre_data[55:48] <= wt_pre_data_w[55:48];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[6] | in_wt_nan[3])) == 1'b0) begin
  end else begin
    wt_pre_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[7] | in_wt_nan[3])) == 1'b1) begin
    wt_pre_data[63:56] <= wt_pre_data_w[63:56];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[7] | in_wt_nan[3])) == 1'b0) begin
  end else begin
    wt_pre_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[8] | in_wt_nan[4])) == 1'b1) begin
    wt_pre_data[71:64] <= wt_pre_data_w[71:64];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[8] | in_wt_nan[4])) == 1'b0) begin
  end else begin
    wt_pre_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[9] | in_wt_nan[4])) == 1'b1) begin
    wt_pre_data[79:72] <= wt_pre_data_w[79:72];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[9] | in_wt_nan[4])) == 1'b0) begin
  end else begin
    wt_pre_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[10] | in_wt_nan[5])) == 1'b1) begin
    wt_pre_data[87:80] <= wt_pre_data_w[87:80];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[10] | in_wt_nan[5])) == 1'b0) begin
  end else begin
    wt_pre_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[11] | in_wt_nan[5])) == 1'b1) begin
    wt_pre_data[95:88] <= wt_pre_data_w[95:88];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[11] | in_wt_nan[5])) == 1'b0) begin
  end else begin
    wt_pre_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[12] | in_wt_nan[6])) == 1'b1) begin
    wt_pre_data[103:96] <= wt_pre_data_w[103:96];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[12] | in_wt_nan[6])) == 1'b0) begin
  end else begin
    wt_pre_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[13] | in_wt_nan[6])) == 1'b1) begin
    wt_pre_data[111:104] <= wt_pre_data_w[111:104];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[13] | in_wt_nan[6])) == 1'b0) begin
  end else begin
    wt_pre_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[14] | in_wt_nan[7])) == 1'b1) begin
    wt_pre_data[119:112] <= wt_pre_data_w[119:112];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[14] | in_wt_nan[7])) == 1'b0) begin
  end else begin
    wt_pre_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[15] | in_wt_nan[7])) == 1'b1) begin
    wt_pre_data[127:120] <= wt_pre_data_w[127:120];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[15] | in_wt_nan[7])) == 1'b0) begin
  end else begin
    wt_pre_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[16] | in_wt_nan[8])) == 1'b1) begin
    wt_pre_data[135:128] <= wt_pre_data_w[135:128];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[16] | in_wt_nan[8])) == 1'b0) begin
  end else begin
    wt_pre_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[17] | in_wt_nan[8])) == 1'b1) begin
    wt_pre_data[143:136] <= wt_pre_data_w[143:136];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[17] | in_wt_nan[8])) == 1'b0) begin
  end else begin
    wt_pre_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[18] | in_wt_nan[9])) == 1'b1) begin
    wt_pre_data[151:144] <= wt_pre_data_w[151:144];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[18] | in_wt_nan[9])) == 1'b0) begin
  end else begin
    wt_pre_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[19] | in_wt_nan[9])) == 1'b1) begin
    wt_pre_data[159:152] <= wt_pre_data_w[159:152];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[19] | in_wt_nan[9])) == 1'b0) begin
  end else begin
    wt_pre_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[20] | in_wt_nan[10])) == 1'b1) begin
    wt_pre_data[167:160] <= wt_pre_data_w[167:160];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[20] | in_wt_nan[10])) == 1'b0) begin
  end else begin
    wt_pre_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[21] | in_wt_nan[10])) == 1'b1) begin
    wt_pre_data[175:168] <= wt_pre_data_w[175:168];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[21] | in_wt_nan[10])) == 1'b0) begin
  end else begin
    wt_pre_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[22] | in_wt_nan[11])) == 1'b1) begin
    wt_pre_data[183:176] <= wt_pre_data_w[183:176];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[22] | in_wt_nan[11])) == 1'b0) begin
  end else begin
    wt_pre_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[23] | in_wt_nan[11])) == 1'b1) begin
    wt_pre_data[191:184] <= wt_pre_data_w[191:184];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[23] | in_wt_nan[11])) == 1'b0) begin
  end else begin
    wt_pre_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[24] | in_wt_nan[12])) == 1'b1) begin
    wt_pre_data[199:192] <= wt_pre_data_w[199:192];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[24] | in_wt_nan[12])) == 1'b0) begin
  end else begin
    wt_pre_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[25] | in_wt_nan[12])) == 1'b1) begin
    wt_pre_data[207:200] <= wt_pre_data_w[207:200];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[25] | in_wt_nan[12])) == 1'b0) begin
  end else begin
    wt_pre_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[26] | in_wt_nan[13])) == 1'b1) begin
    wt_pre_data[215:208] <= wt_pre_data_w[215:208];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[26] | in_wt_nan[13])) == 1'b0) begin
  end else begin
    wt_pre_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[27] | in_wt_nan[13])) == 1'b1) begin
    wt_pre_data[223:216] <= wt_pre_data_w[223:216];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[27] | in_wt_nan[13])) == 1'b0) begin
  end else begin
    wt_pre_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[28] | in_wt_nan[14])) == 1'b1) begin
    wt_pre_data[231:224] <= wt_pre_data_w[231:224];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[28] | in_wt_nan[14])) == 1'b0) begin
  end else begin
    wt_pre_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[29] | in_wt_nan[14])) == 1'b1) begin
    wt_pre_data[239:232] <= wt_pre_data_w[239:232];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[29] | in_wt_nan[14])) == 1'b0) begin
  end else begin
    wt_pre_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[30] | in_wt_nan[15])) == 1'b1) begin
    wt_pre_data[247:240] <= wt_pre_data_w[247:240];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[30] | in_wt_nan[15])) == 1'b0) begin
  end else begin
    wt_pre_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[31] | in_wt_nan[15])) == 1'b1) begin
    wt_pre_data[255:248] <= wt_pre_data_w[255:248];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[31] | in_wt_nan[15])) == 1'b0) begin
  end else begin
    wt_pre_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[32] | in_wt_nan[16])) == 1'b1) begin
    wt_pre_data[263:256] <= wt_pre_data_w[263:256];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[32] | in_wt_nan[16])) == 1'b0) begin
  end else begin
    wt_pre_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[33] | in_wt_nan[16])) == 1'b1) begin
    wt_pre_data[271:264] <= wt_pre_data_w[271:264];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[33] | in_wt_nan[16])) == 1'b0) begin
  end else begin
    wt_pre_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[34] | in_wt_nan[17])) == 1'b1) begin
    wt_pre_data[279:272] <= wt_pre_data_w[279:272];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[34] | in_wt_nan[17])) == 1'b0) begin
  end else begin
    wt_pre_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[35] | in_wt_nan[17])) == 1'b1) begin
    wt_pre_data[287:280] <= wt_pre_data_w[287:280];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[35] | in_wt_nan[17])) == 1'b0) begin
  end else begin
    wt_pre_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[36] | in_wt_nan[18])) == 1'b1) begin
    wt_pre_data[295:288] <= wt_pre_data_w[295:288];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[36] | in_wt_nan[18])) == 1'b0) begin
  end else begin
    wt_pre_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[37] | in_wt_nan[18])) == 1'b1) begin
    wt_pre_data[303:296] <= wt_pre_data_w[303:296];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[37] | in_wt_nan[18])) == 1'b0) begin
  end else begin
    wt_pre_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[38] | in_wt_nan[19])) == 1'b1) begin
    wt_pre_data[311:304] <= wt_pre_data_w[311:304];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[38] | in_wt_nan[19])) == 1'b0) begin
  end else begin
    wt_pre_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[39] | in_wt_nan[19])) == 1'b1) begin
    wt_pre_data[319:312] <= wt_pre_data_w[319:312];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[39] | in_wt_nan[19])) == 1'b0) begin
  end else begin
    wt_pre_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[40] | in_wt_nan[20])) == 1'b1) begin
    wt_pre_data[327:320] <= wt_pre_data_w[327:320];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[40] | in_wt_nan[20])) == 1'b0) begin
  end else begin
    wt_pre_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[41] | in_wt_nan[20])) == 1'b1) begin
    wt_pre_data[335:328] <= wt_pre_data_w[335:328];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[41] | in_wt_nan[20])) == 1'b0) begin
  end else begin
    wt_pre_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[42] | in_wt_nan[21])) == 1'b1) begin
    wt_pre_data[343:336] <= wt_pre_data_w[343:336];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[42] | in_wt_nan[21])) == 1'b0) begin
  end else begin
    wt_pre_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[43] | in_wt_nan[21])) == 1'b1) begin
    wt_pre_data[351:344] <= wt_pre_data_w[351:344];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[43] | in_wt_nan[21])) == 1'b0) begin
  end else begin
    wt_pre_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[44] | in_wt_nan[22])) == 1'b1) begin
    wt_pre_data[359:352] <= wt_pre_data_w[359:352];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[44] | in_wt_nan[22])) == 1'b0) begin
  end else begin
    wt_pre_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[45] | in_wt_nan[22])) == 1'b1) begin
    wt_pre_data[367:360] <= wt_pre_data_w[367:360];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[45] | in_wt_nan[22])) == 1'b0) begin
  end else begin
    wt_pre_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[46] | in_wt_nan[23])) == 1'b1) begin
    wt_pre_data[375:368] <= wt_pre_data_w[375:368];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[46] | in_wt_nan[23])) == 1'b0) begin
  end else begin
    wt_pre_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[47] | in_wt_nan[23])) == 1'b1) begin
    wt_pre_data[383:376] <= wt_pre_data_w[383:376];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[47] | in_wt_nan[23])) == 1'b0) begin
  end else begin
    wt_pre_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[48] | in_wt_nan[24])) == 1'b1) begin
    wt_pre_data[391:384] <= wt_pre_data_w[391:384];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[48] | in_wt_nan[24])) == 1'b0) begin
  end else begin
    wt_pre_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[49] | in_wt_nan[24])) == 1'b1) begin
    wt_pre_data[399:392] <= wt_pre_data_w[399:392];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[49] | in_wt_nan[24])) == 1'b0) begin
  end else begin
    wt_pre_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[50] | in_wt_nan[25])) == 1'b1) begin
    wt_pre_data[407:400] <= wt_pre_data_w[407:400];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[50] | in_wt_nan[25])) == 1'b0) begin
  end else begin
    wt_pre_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[51] | in_wt_nan[25])) == 1'b1) begin
    wt_pre_data[415:408] <= wt_pre_data_w[415:408];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[51] | in_wt_nan[25])) == 1'b0) begin
  end else begin
    wt_pre_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[52] | in_wt_nan[26])) == 1'b1) begin
    wt_pre_data[423:416] <= wt_pre_data_w[423:416];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[52] | in_wt_nan[26])) == 1'b0) begin
  end else begin
    wt_pre_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[53] | in_wt_nan[26])) == 1'b1) begin
    wt_pre_data[431:424] <= wt_pre_data_w[431:424];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[53] | in_wt_nan[26])) == 1'b0) begin
  end else begin
    wt_pre_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[54] | in_wt_nan[27])) == 1'b1) begin
    wt_pre_data[439:432] <= wt_pre_data_w[439:432];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[54] | in_wt_nan[27])) == 1'b0) begin
  end else begin
    wt_pre_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[55] | in_wt_nan[27])) == 1'b1) begin
    wt_pre_data[447:440] <= wt_pre_data_w[447:440];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[55] | in_wt_nan[27])) == 1'b0) begin
  end else begin
    wt_pre_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[56] | in_wt_nan[28])) == 1'b1) begin
    wt_pre_data[455:448] <= wt_pre_data_w[455:448];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[56] | in_wt_nan[28])) == 1'b0) begin
  end else begin
    wt_pre_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[57] | in_wt_nan[28])) == 1'b1) begin
    wt_pre_data[463:456] <= wt_pre_data_w[463:456];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[57] | in_wt_nan[28])) == 1'b0) begin
  end else begin
    wt_pre_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[58] | in_wt_nan[29])) == 1'b1) begin
    wt_pre_data[471:464] <= wt_pre_data_w[471:464];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[58] | in_wt_nan[29])) == 1'b0) begin
  end else begin
    wt_pre_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[59] | in_wt_nan[29])) == 1'b1) begin
    wt_pre_data[479:472] <= wt_pre_data_w[479:472];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[59] | in_wt_nan[29])) == 1'b0) begin
  end else begin
    wt_pre_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[60] | in_wt_nan[30])) == 1'b1) begin
    wt_pre_data[487:480] <= wt_pre_data_w[487:480];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[60] | in_wt_nan[30])) == 1'b0) begin
  end else begin
    wt_pre_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[61] | in_wt_nan[30])) == 1'b1) begin
    wt_pre_data[495:488] <= wt_pre_data_w[495:488];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[61] | in_wt_nan[30])) == 1'b0) begin
  end else begin
    wt_pre_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[62] | in_wt_nan[31])) == 1'b1) begin
    wt_pre_data[503:496] <= wt_pre_data_w[503:496];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[62] | in_wt_nan[31])) == 1'b0) begin
  end else begin
    wt_pre_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[63] | in_wt_nan[31])) == 1'b1) begin
    wt_pre_data[511:504] <= wt_pre_data_w[511:504];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[63] | in_wt_nan[31])) == 1'b0) begin
  end else begin
    wt_pre_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[64] | in_wt_nan[32])) == 1'b1) begin
    wt_pre_data[519:512] <= wt_pre_data_w[519:512];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[64] | in_wt_nan[32])) == 1'b0) begin
  end else begin
    wt_pre_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[65] | in_wt_nan[32])) == 1'b1) begin
    wt_pre_data[527:520] <= wt_pre_data_w[527:520];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[65] | in_wt_nan[32])) == 1'b0) begin
  end else begin
    wt_pre_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[66] | in_wt_nan[33])) == 1'b1) begin
    wt_pre_data[535:528] <= wt_pre_data_w[535:528];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[66] | in_wt_nan[33])) == 1'b0) begin
  end else begin
    wt_pre_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[67] | in_wt_nan[33])) == 1'b1) begin
    wt_pre_data[543:536] <= wt_pre_data_w[543:536];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[67] | in_wt_nan[33])) == 1'b0) begin
  end else begin
    wt_pre_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[68] | in_wt_nan[34])) == 1'b1) begin
    wt_pre_data[551:544] <= wt_pre_data_w[551:544];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[68] | in_wt_nan[34])) == 1'b0) begin
  end else begin
    wt_pre_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[69] | in_wt_nan[34])) == 1'b1) begin
    wt_pre_data[559:552] <= wt_pre_data_w[559:552];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[69] | in_wt_nan[34])) == 1'b0) begin
  end else begin
    wt_pre_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[70] | in_wt_nan[35])) == 1'b1) begin
    wt_pre_data[567:560] <= wt_pre_data_w[567:560];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[70] | in_wt_nan[35])) == 1'b0) begin
  end else begin
    wt_pre_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[71] | in_wt_nan[35])) == 1'b1) begin
    wt_pre_data[575:568] <= wt_pre_data_w[575:568];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[71] | in_wt_nan[35])) == 1'b0) begin
  end else begin
    wt_pre_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[72] | in_wt_nan[36])) == 1'b1) begin
    wt_pre_data[583:576] <= wt_pre_data_w[583:576];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[72] | in_wt_nan[36])) == 1'b0) begin
  end else begin
    wt_pre_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[73] | in_wt_nan[36])) == 1'b1) begin
    wt_pre_data[591:584] <= wt_pre_data_w[591:584];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[73] | in_wt_nan[36])) == 1'b0) begin
  end else begin
    wt_pre_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[74] | in_wt_nan[37])) == 1'b1) begin
    wt_pre_data[599:592] <= wt_pre_data_w[599:592];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[74] | in_wt_nan[37])) == 1'b0) begin
  end else begin
    wt_pre_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[75] | in_wt_nan[37])) == 1'b1) begin
    wt_pre_data[607:600] <= wt_pre_data_w[607:600];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[75] | in_wt_nan[37])) == 1'b0) begin
  end else begin
    wt_pre_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[76] | in_wt_nan[38])) == 1'b1) begin
    wt_pre_data[615:608] <= wt_pre_data_w[615:608];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[76] | in_wt_nan[38])) == 1'b0) begin
  end else begin
    wt_pre_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[77] | in_wt_nan[38])) == 1'b1) begin
    wt_pre_data[623:616] <= wt_pre_data_w[623:616];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[77] | in_wt_nan[38])) == 1'b0) begin
  end else begin
    wt_pre_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[78] | in_wt_nan[39])) == 1'b1) begin
    wt_pre_data[631:624] <= wt_pre_data_w[631:624];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[78] | in_wt_nan[39])) == 1'b0) begin
  end else begin
    wt_pre_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[79] | in_wt_nan[39])) == 1'b1) begin
    wt_pre_data[639:632] <= wt_pre_data_w[639:632];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[79] | in_wt_nan[39])) == 1'b0) begin
  end else begin
    wt_pre_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[80] | in_wt_nan[40])) == 1'b1) begin
    wt_pre_data[647:640] <= wt_pre_data_w[647:640];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[80] | in_wt_nan[40])) == 1'b0) begin
  end else begin
    wt_pre_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[81] | in_wt_nan[40])) == 1'b1) begin
    wt_pre_data[655:648] <= wt_pre_data_w[655:648];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[81] | in_wt_nan[40])) == 1'b0) begin
  end else begin
    wt_pre_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[82] | in_wt_nan[41])) == 1'b1) begin
    wt_pre_data[663:656] <= wt_pre_data_w[663:656];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[82] | in_wt_nan[41])) == 1'b0) begin
  end else begin
    wt_pre_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[83] | in_wt_nan[41])) == 1'b1) begin
    wt_pre_data[671:664] <= wt_pre_data_w[671:664];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[83] | in_wt_nan[41])) == 1'b0) begin
  end else begin
    wt_pre_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[84] | in_wt_nan[42])) == 1'b1) begin
    wt_pre_data[679:672] <= wt_pre_data_w[679:672];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[84] | in_wt_nan[42])) == 1'b0) begin
  end else begin
    wt_pre_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[85] | in_wt_nan[42])) == 1'b1) begin
    wt_pre_data[687:680] <= wt_pre_data_w[687:680];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[85] | in_wt_nan[42])) == 1'b0) begin
  end else begin
    wt_pre_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[86] | in_wt_nan[43])) == 1'b1) begin
    wt_pre_data[695:688] <= wt_pre_data_w[695:688];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[86] | in_wt_nan[43])) == 1'b0) begin
  end else begin
    wt_pre_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[87] | in_wt_nan[43])) == 1'b1) begin
    wt_pre_data[703:696] <= wt_pre_data_w[703:696];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[87] | in_wt_nan[43])) == 1'b0) begin
  end else begin
    wt_pre_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[88] | in_wt_nan[44])) == 1'b1) begin
    wt_pre_data[711:704] <= wt_pre_data_w[711:704];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[88] | in_wt_nan[44])) == 1'b0) begin
  end else begin
    wt_pre_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[89] | in_wt_nan[44])) == 1'b1) begin
    wt_pre_data[719:712] <= wt_pre_data_w[719:712];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[89] | in_wt_nan[44])) == 1'b0) begin
  end else begin
    wt_pre_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[90] | in_wt_nan[45])) == 1'b1) begin
    wt_pre_data[727:720] <= wt_pre_data_w[727:720];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[90] | in_wt_nan[45])) == 1'b0) begin
  end else begin
    wt_pre_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[91] | in_wt_nan[45])) == 1'b1) begin
    wt_pre_data[735:728] <= wt_pre_data_w[735:728];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[91] | in_wt_nan[45])) == 1'b0) begin
  end else begin
    wt_pre_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[92] | in_wt_nan[46])) == 1'b1) begin
    wt_pre_data[743:736] <= wt_pre_data_w[743:736];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[92] | in_wt_nan[46])) == 1'b0) begin
  end else begin
    wt_pre_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[93] | in_wt_nan[46])) == 1'b1) begin
    wt_pre_data[751:744] <= wt_pre_data_w[751:744];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[93] | in_wt_nan[46])) == 1'b0) begin
  end else begin
    wt_pre_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[94] | in_wt_nan[47])) == 1'b1) begin
    wt_pre_data[759:752] <= wt_pre_data_w[759:752];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[94] | in_wt_nan[47])) == 1'b0) begin
  end else begin
    wt_pre_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[95] | in_wt_nan[47])) == 1'b1) begin
    wt_pre_data[767:760] <= wt_pre_data_w[767:760];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[95] | in_wt_nan[47])) == 1'b0) begin
  end else begin
    wt_pre_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[96] | in_wt_nan[48])) == 1'b1) begin
    wt_pre_data[775:768] <= wt_pre_data_w[775:768];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[96] | in_wt_nan[48])) == 1'b0) begin
  end else begin
    wt_pre_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[97] | in_wt_nan[48])) == 1'b1) begin
    wt_pre_data[783:776] <= wt_pre_data_w[783:776];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[97] | in_wt_nan[48])) == 1'b0) begin
  end else begin
    wt_pre_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[98] | in_wt_nan[49])) == 1'b1) begin
    wt_pre_data[791:784] <= wt_pre_data_w[791:784];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[98] | in_wt_nan[49])) == 1'b0) begin
  end else begin
    wt_pre_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[99] | in_wt_nan[49])) == 1'b1) begin
    wt_pre_data[799:792] <= wt_pre_data_w[799:792];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[99] | in_wt_nan[49])) == 1'b0) begin
  end else begin
    wt_pre_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[100] | in_wt_nan[50])) == 1'b1) begin
    wt_pre_data[807:800] <= wt_pre_data_w[807:800];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[100] | in_wt_nan[50])) == 1'b0) begin
  end else begin
    wt_pre_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[101] | in_wt_nan[50])) == 1'b1) begin
    wt_pre_data[815:808] <= wt_pre_data_w[815:808];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[101] | in_wt_nan[50])) == 1'b0) begin
  end else begin
    wt_pre_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[102] | in_wt_nan[51])) == 1'b1) begin
    wt_pre_data[823:816] <= wt_pre_data_w[823:816];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[102] | in_wt_nan[51])) == 1'b0) begin
  end else begin
    wt_pre_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[103] | in_wt_nan[51])) == 1'b1) begin
    wt_pre_data[831:824] <= wt_pre_data_w[831:824];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[103] | in_wt_nan[51])) == 1'b0) begin
  end else begin
    wt_pre_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[104] | in_wt_nan[52])) == 1'b1) begin
    wt_pre_data[839:832] <= wt_pre_data_w[839:832];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[104] | in_wt_nan[52])) == 1'b0) begin
  end else begin
    wt_pre_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[105] | in_wt_nan[52])) == 1'b1) begin
    wt_pre_data[847:840] <= wt_pre_data_w[847:840];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[105] | in_wt_nan[52])) == 1'b0) begin
  end else begin
    wt_pre_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[106] | in_wt_nan[53])) == 1'b1) begin
    wt_pre_data[855:848] <= wt_pre_data_w[855:848];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[106] | in_wt_nan[53])) == 1'b0) begin
  end else begin
    wt_pre_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[107] | in_wt_nan[53])) == 1'b1) begin
    wt_pre_data[863:856] <= wt_pre_data_w[863:856];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[107] | in_wt_nan[53])) == 1'b0) begin
  end else begin
    wt_pre_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[108] | in_wt_nan[54])) == 1'b1) begin
    wt_pre_data[871:864] <= wt_pre_data_w[871:864];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[108] | in_wt_nan[54])) == 1'b0) begin
  end else begin
    wt_pre_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[109] | in_wt_nan[54])) == 1'b1) begin
    wt_pre_data[879:872] <= wt_pre_data_w[879:872];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[109] | in_wt_nan[54])) == 1'b0) begin
  end else begin
    wt_pre_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[110] | in_wt_nan[55])) == 1'b1) begin
    wt_pre_data[887:880] <= wt_pre_data_w[887:880];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[110] | in_wt_nan[55])) == 1'b0) begin
  end else begin
    wt_pre_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[111] | in_wt_nan[55])) == 1'b1) begin
    wt_pre_data[895:888] <= wt_pre_data_w[895:888];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[111] | in_wt_nan[55])) == 1'b0) begin
  end else begin
    wt_pre_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[112] | in_wt_nan[56])) == 1'b1) begin
    wt_pre_data[903:896] <= wt_pre_data_w[903:896];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[112] | in_wt_nan[56])) == 1'b0) begin
  end else begin
    wt_pre_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[113] | in_wt_nan[56])) == 1'b1) begin
    wt_pre_data[911:904] <= wt_pre_data_w[911:904];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[113] | in_wt_nan[56])) == 1'b0) begin
  end else begin
    wt_pre_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[114] | in_wt_nan[57])) == 1'b1) begin
    wt_pre_data[919:912] <= wt_pre_data_w[919:912];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[114] | in_wt_nan[57])) == 1'b0) begin
  end else begin
    wt_pre_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[115] | in_wt_nan[57])) == 1'b1) begin
    wt_pre_data[927:920] <= wt_pre_data_w[927:920];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[115] | in_wt_nan[57])) == 1'b0) begin
  end else begin
    wt_pre_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[116] | in_wt_nan[58])) == 1'b1) begin
    wt_pre_data[935:928] <= wt_pre_data_w[935:928];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[116] | in_wt_nan[58])) == 1'b0) begin
  end else begin
    wt_pre_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[117] | in_wt_nan[58])) == 1'b1) begin
    wt_pre_data[943:936] <= wt_pre_data_w[943:936];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[117] | in_wt_nan[58])) == 1'b0) begin
  end else begin
    wt_pre_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[118] | in_wt_nan[59])) == 1'b1) begin
    wt_pre_data[951:944] <= wt_pre_data_w[951:944];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[118] | in_wt_nan[59])) == 1'b0) begin
  end else begin
    wt_pre_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[119] | in_wt_nan[59])) == 1'b1) begin
    wt_pre_data[959:952] <= wt_pre_data_w[959:952];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[119] | in_wt_nan[59])) == 1'b0) begin
  end else begin
    wt_pre_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[120] | in_wt_nan[60])) == 1'b1) begin
    wt_pre_data[967:960] <= wt_pre_data_w[967:960];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[120] | in_wt_nan[60])) == 1'b0) begin
  end else begin
    wt_pre_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[121] | in_wt_nan[60])) == 1'b1) begin
    wt_pre_data[975:968] <= wt_pre_data_w[975:968];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[121] | in_wt_nan[60])) == 1'b0) begin
  end else begin
    wt_pre_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[122] | in_wt_nan[61])) == 1'b1) begin
    wt_pre_data[983:976] <= wt_pre_data_w[983:976];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[122] | in_wt_nan[61])) == 1'b0) begin
  end else begin
    wt_pre_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[123] | in_wt_nan[61])) == 1'b1) begin
    wt_pre_data[991:984] <= wt_pre_data_w[991:984];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[123] | in_wt_nan[61])) == 1'b0) begin
  end else begin
    wt_pre_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[124] | in_wt_nan[62])) == 1'b1) begin
    wt_pre_data[999:992] <= wt_pre_data_w[999:992];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[124] | in_wt_nan[62])) == 1'b0) begin
  end else begin
    wt_pre_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[125] | in_wt_nan[62])) == 1'b1) begin
    wt_pre_data[1007:1000] <= wt_pre_data_w[1007:1000];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[125] | in_wt_nan[62])) == 1'b0) begin
  end else begin
    wt_pre_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[126] | in_wt_nan[63])) == 1'b1) begin
    wt_pre_data[1015:1008] <= wt_pre_data_w[1015:1008];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[126] | in_wt_nan[63])) == 1'b0) begin
  end else begin
    wt_pre_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_wt_pvld & (wt_pre_nz_w[127] | in_wt_nan[63])) == 1'b1) begin
    wt_pre_data[1023:1016] <= wt_pre_data_w[1023:1016];
  // VCS coverage off
  end else if ((in_wt_pvld & (wt_pre_nz_w[127] | in_wt_nan[63])) == 1'b0) begin
  end else begin
    wt_pre_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

//==========================================================
// Weight shawdow and active register         
//==========================================================


always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt0_sd_pvld
  ) begin
    wt0_sd_pvld_w = wt_pre_sel[0] ? 1'b1 :
                    dat_pre_stripe_st[0] ? 1'b0 :
                    wt0_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt0_sd_pvld <= 1'b0;
  end else begin
  wt0_sd_pvld <= wt0_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0]) == 1'b1) begin
    wt0_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[0]) == 1'b0) begin
  end else begin
    wt0_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b1) begin
    wt0_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b0) begin
  end else begin
    wt0_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b1) begin
    wt0_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b0) begin
  end else begin
    wt0_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b1) begin
    wt0_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[0] & cfg_is_fp16_d1[66]) == 1'b0) begin
  end else begin
    wt0_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt0_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt0_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt0_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt0_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt0_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt0_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt0_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt0_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt0_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt0_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt0_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt0_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt0_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt0_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt0_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt0_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt0_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt0_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt0_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt0_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt0_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt0_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt0_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt0_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt0_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt0_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt0_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt0_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt0_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt0_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt0_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt0_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt0_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt0_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt0_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt0_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt0_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt0_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt0_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt0_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt0_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt0_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt0_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt0_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt0_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt0_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt0_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt0_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt0_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt0_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt0_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt0_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt0_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt0_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt0_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt0_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt0_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt0_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt0_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt0_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt0_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt0_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt0_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt0_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt0_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt0_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt0_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt0_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt0_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt0_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt0_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt0_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt0_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt0_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt0_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt0_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt0_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt0_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt0_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt0_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt0_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt0_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt0_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt0_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt0_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt0_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt0_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt0_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt0_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt0_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt0_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt0_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt0_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt0_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt0_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt0_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt0_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt0_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt0_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt0_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt0_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt0_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt0_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt0_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt0_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt0_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt0_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt0_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt0_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt0_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt0_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt0_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt0_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt0_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt0_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt0_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt0_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt0_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt0_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt0_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt0_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt0_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt0_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt0_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt0_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt0_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt0_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt0_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt0_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt0_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt0_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt0_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt0_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt0_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt0_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt0_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt0_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt0_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt0_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt0_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt0_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt0_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt0_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt0_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt0_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt0_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt0_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt0_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt0_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt0_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt0_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt0_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt0_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt0_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt0_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt0_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt0_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt0_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt0_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt0_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt0_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt0_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt0_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt0_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt0_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt0_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt0_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt0_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt0_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt0_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt0_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt0_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt0_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt0_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt0_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt0_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt0_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt0_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt0_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt0_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt0_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt0_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt0_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt0_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt0_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt0_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt0_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt0_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt0_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt0_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt0_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt0_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt0_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt0_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt0_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt0_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt0_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt0_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt0_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt0_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt0_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt0_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt0_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt0_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt0_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt0_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt0_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt0_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt0_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt0_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt0_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt0_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt0_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt0_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt0_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt0_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt0_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt0_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt0_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt0_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt0_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt0_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt0_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt0_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt0_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt0_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt0_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt0_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt0_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt0_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt0_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt0_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt0_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt0_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt0_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt0_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt0_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt0_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt0_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt0_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt0_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt0_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt0_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt0_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt0_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt0_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt0_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt0_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt0_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt0_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt0_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt0_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt0_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt0_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[0] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt0_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[0] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt0_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt1_sd_pvld
  ) begin
    wt1_sd_pvld_w = wt_pre_sel[1] ? 1'b1 :
                    dat_pre_stripe_st[1] ? 1'b0 :
                    wt1_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt1_sd_pvld <= 1'b0;
  end else begin
  wt1_sd_pvld <= wt1_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1]) == 1'b1) begin
    wt1_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[1]) == 1'b0) begin
  end else begin
    wt1_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b1) begin
    wt1_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b0) begin
  end else begin
    wt1_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b1) begin
    wt1_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b0) begin
  end else begin
    wt1_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b1) begin
    wt1_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[1] & cfg_is_fp16_d1[67]) == 1'b0) begin
  end else begin
    wt1_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt1_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt1_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt1_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt1_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt1_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt1_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt1_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt1_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt1_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt1_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt1_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt1_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt1_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt1_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt1_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt1_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt1_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt1_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt1_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt1_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt1_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt1_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt1_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt1_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt1_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt1_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt1_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt1_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt1_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt1_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt1_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt1_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt1_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt1_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt1_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt1_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt1_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt1_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt1_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt1_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt1_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt1_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt1_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt1_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt1_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt1_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt1_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt1_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt1_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt1_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt1_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt1_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt1_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt1_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt1_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt1_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt1_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt1_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt1_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt1_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt1_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt1_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt1_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt1_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt1_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt1_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt1_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt1_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt1_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt1_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt1_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt1_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt1_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt1_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt1_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt1_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt1_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt1_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt1_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt1_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt1_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt1_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt1_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt1_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt1_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt1_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt1_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt1_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt1_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt1_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt1_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt1_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt1_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt1_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt1_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt1_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt1_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt1_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt1_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt1_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt1_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt1_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt1_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt1_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt1_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt1_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt1_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt1_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt1_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt1_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt1_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt1_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt1_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt1_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt1_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt1_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt1_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt1_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt1_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt1_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt1_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt1_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt1_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt1_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt1_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt1_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt1_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt1_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt1_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt1_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt1_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt1_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt1_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt1_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt1_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt1_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt1_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt1_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt1_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt1_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt1_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt1_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt1_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt1_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt1_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt1_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt1_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt1_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt1_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt1_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt1_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt1_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt1_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt1_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt1_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt1_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt1_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt1_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt1_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt1_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt1_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt1_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt1_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt1_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt1_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt1_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt1_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt1_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt1_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt1_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt1_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt1_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt1_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt1_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt1_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt1_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt1_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt1_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt1_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt1_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt1_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt1_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt1_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt1_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt1_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt1_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt1_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt1_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt1_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt1_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt1_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt1_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt1_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt1_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt1_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt1_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt1_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt1_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt1_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt1_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt1_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt1_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt1_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt1_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt1_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt1_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt1_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt1_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt1_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt1_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt1_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt1_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt1_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt1_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt1_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt1_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt1_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt1_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt1_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt1_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt1_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt1_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt1_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt1_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt1_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt1_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt1_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt1_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt1_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt1_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt1_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt1_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt1_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt1_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt1_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt1_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt1_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt1_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt1_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt1_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt1_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt1_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt1_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt1_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt1_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt1_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt1_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt1_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt1_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt1_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt1_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt1_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt1_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt1_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[1] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt1_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[1] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt1_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt2_sd_pvld
  ) begin
    wt2_sd_pvld_w = wt_pre_sel[2] ? 1'b1 :
                    dat_pre_stripe_st[2] ? 1'b0 :
                    wt2_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt2_sd_pvld <= 1'b0;
  end else begin
  wt2_sd_pvld <= wt2_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2]) == 1'b1) begin
    wt2_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[2]) == 1'b0) begin
  end else begin
    wt2_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b1) begin
    wt2_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b0) begin
  end else begin
    wt2_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b1) begin
    wt2_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b0) begin
  end else begin
    wt2_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b1) begin
    wt2_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[2] & cfg_is_fp16_d1[68]) == 1'b0) begin
  end else begin
    wt2_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt2_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt2_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt2_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt2_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt2_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt2_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt2_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt2_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt2_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt2_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt2_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt2_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt2_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt2_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt2_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt2_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt2_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt2_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt2_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt2_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt2_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt2_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt2_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt2_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt2_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt2_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt2_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt2_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt2_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt2_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt2_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt2_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt2_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt2_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt2_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt2_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt2_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt2_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt2_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt2_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt2_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt2_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt2_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt2_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt2_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt2_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt2_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt2_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt2_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt2_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt2_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt2_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt2_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt2_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt2_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt2_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt2_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt2_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt2_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt2_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt2_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt2_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt2_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt2_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt2_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt2_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt2_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt2_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt2_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt2_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt2_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt2_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt2_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt2_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt2_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt2_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt2_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt2_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt2_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt2_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt2_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt2_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt2_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt2_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt2_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt2_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt2_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt2_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt2_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt2_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt2_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt2_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt2_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt2_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt2_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt2_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt2_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt2_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt2_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt2_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt2_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt2_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt2_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt2_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt2_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt2_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt2_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt2_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt2_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt2_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt2_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt2_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt2_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt2_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt2_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt2_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt2_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt2_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt2_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt2_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt2_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt2_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt2_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt2_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt2_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt2_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt2_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt2_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt2_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt2_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt2_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt2_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt2_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt2_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt2_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt2_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt2_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt2_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt2_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt2_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt2_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt2_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt2_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt2_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt2_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt2_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt2_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt2_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt2_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt2_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt2_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt2_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt2_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt2_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt2_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt2_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt2_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt2_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt2_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt2_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt2_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt2_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt2_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt2_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt2_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt2_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt2_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt2_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt2_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt2_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt2_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt2_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt2_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt2_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt2_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt2_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt2_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt2_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt2_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt2_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt2_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt2_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt2_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt2_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt2_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt2_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt2_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt2_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt2_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt2_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt2_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt2_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt2_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt2_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt2_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt2_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt2_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt2_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt2_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt2_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt2_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt2_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt2_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt2_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt2_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt2_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt2_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt2_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt2_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt2_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt2_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt2_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt2_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt2_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt2_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt2_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt2_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt2_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt2_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt2_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt2_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt2_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt2_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt2_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt2_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt2_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt2_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt2_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt2_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt2_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt2_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt2_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt2_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt2_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt2_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt2_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt2_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt2_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt2_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt2_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt2_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt2_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt2_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt2_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt2_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt2_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt2_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt2_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt2_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt2_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt2_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt2_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt2_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt2_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[2] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt2_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[2] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt2_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt3_sd_pvld
  ) begin
    wt3_sd_pvld_w = wt_pre_sel[3] ? 1'b1 :
                    dat_pre_stripe_st[3] ? 1'b0 :
                    wt3_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt3_sd_pvld <= 1'b0;
  end else begin
  wt3_sd_pvld <= wt3_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3]) == 1'b1) begin
    wt3_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[3]) == 1'b0) begin
  end else begin
    wt3_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b1) begin
    wt3_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b0) begin
  end else begin
    wt3_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b1) begin
    wt3_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b0) begin
  end else begin
    wt3_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b1) begin
    wt3_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[3] & cfg_is_fp16_d1[69]) == 1'b0) begin
  end else begin
    wt3_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt3_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt3_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt3_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt3_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt3_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt3_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt3_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt3_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt3_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt3_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt3_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt3_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt3_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt3_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt3_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt3_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt3_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt3_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt3_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt3_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt3_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt3_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt3_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt3_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt3_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt3_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt3_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt3_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt3_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt3_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt3_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt3_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt3_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt3_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt3_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt3_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt3_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt3_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt3_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt3_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt3_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt3_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt3_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt3_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt3_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt3_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt3_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt3_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt3_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt3_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt3_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt3_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt3_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt3_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt3_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt3_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt3_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt3_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt3_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt3_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt3_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt3_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt3_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt3_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt3_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt3_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt3_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt3_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt3_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt3_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt3_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt3_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt3_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt3_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt3_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt3_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt3_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt3_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt3_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt3_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt3_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt3_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt3_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt3_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt3_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt3_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt3_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt3_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt3_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt3_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt3_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt3_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt3_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt3_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt3_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt3_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt3_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt3_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt3_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt3_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt3_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt3_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt3_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt3_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt3_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt3_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt3_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt3_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt3_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt3_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt3_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt3_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt3_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt3_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt3_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt3_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt3_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt3_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt3_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt3_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt3_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt3_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt3_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt3_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt3_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt3_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt3_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt3_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt3_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt3_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt3_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt3_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt3_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt3_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt3_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt3_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt3_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt3_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt3_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt3_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt3_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt3_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt3_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt3_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt3_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt3_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt3_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt3_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt3_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt3_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt3_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt3_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt3_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt3_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt3_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt3_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt3_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt3_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt3_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt3_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt3_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt3_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt3_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt3_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt3_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt3_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt3_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt3_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt3_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt3_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt3_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt3_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt3_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt3_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt3_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt3_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt3_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt3_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt3_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt3_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt3_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt3_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt3_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt3_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt3_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt3_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt3_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt3_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt3_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt3_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt3_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt3_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt3_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt3_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt3_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt3_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt3_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt3_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt3_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt3_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt3_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt3_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt3_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt3_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt3_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt3_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt3_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt3_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt3_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt3_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt3_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt3_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt3_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt3_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt3_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt3_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt3_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt3_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt3_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt3_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt3_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt3_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt3_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt3_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt3_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt3_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt3_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt3_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt3_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt3_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt3_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt3_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt3_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt3_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt3_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt3_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt3_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt3_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt3_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt3_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt3_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt3_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt3_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt3_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt3_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt3_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt3_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt3_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt3_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt3_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt3_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt3_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt3_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt3_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[3] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt3_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[3] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt3_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt4_sd_pvld
  ) begin
    wt4_sd_pvld_w = wt_pre_sel[4] ? 1'b1 :
                    dat_pre_stripe_st[4] ? 1'b0 :
                    wt4_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt4_sd_pvld <= 1'b0;
  end else begin
  wt4_sd_pvld <= wt4_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4]) == 1'b1) begin
    wt4_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[4]) == 1'b0) begin
  end else begin
    wt4_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b1) begin
    wt4_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b0) begin
  end else begin
    wt4_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b1) begin
    wt4_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b0) begin
  end else begin
    wt4_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b1) begin
    wt4_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[4] & cfg_is_fp16_d1[70]) == 1'b0) begin
  end else begin
    wt4_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt4_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt4_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt4_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt4_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt4_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt4_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt4_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt4_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt4_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt4_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt4_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt4_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt4_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt4_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt4_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt4_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt4_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt4_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt4_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt4_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt4_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt4_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt4_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt4_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt4_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt4_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt4_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt4_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt4_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt4_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt4_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt4_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt4_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt4_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt4_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt4_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt4_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt4_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt4_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt4_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt4_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt4_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt4_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt4_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt4_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt4_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt4_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt4_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt4_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt4_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt4_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt4_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt4_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt4_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt4_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt4_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt4_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt4_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt4_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt4_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt4_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt4_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt4_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt4_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt4_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt4_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt4_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt4_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt4_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt4_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt4_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt4_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt4_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt4_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt4_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt4_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt4_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt4_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt4_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt4_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt4_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt4_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt4_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt4_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt4_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt4_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt4_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt4_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt4_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt4_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt4_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt4_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt4_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt4_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt4_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt4_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt4_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt4_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt4_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt4_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt4_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt4_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt4_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt4_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt4_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt4_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt4_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt4_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt4_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt4_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt4_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt4_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt4_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt4_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt4_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt4_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt4_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt4_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt4_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt4_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt4_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt4_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt4_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt4_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt4_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt4_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt4_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt4_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt4_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt4_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt4_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt4_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt4_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt4_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt4_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt4_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt4_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt4_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt4_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt4_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt4_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt4_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt4_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt4_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt4_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt4_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt4_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt4_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt4_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt4_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt4_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt4_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt4_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt4_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt4_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt4_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt4_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt4_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt4_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt4_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt4_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt4_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt4_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt4_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt4_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt4_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt4_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt4_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt4_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt4_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt4_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt4_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt4_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt4_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt4_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt4_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt4_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt4_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt4_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt4_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt4_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt4_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt4_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt4_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt4_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt4_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt4_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt4_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt4_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt4_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt4_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt4_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt4_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt4_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt4_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt4_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt4_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt4_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt4_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt4_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt4_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt4_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt4_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt4_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt4_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt4_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt4_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt4_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt4_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt4_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt4_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt4_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt4_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt4_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt4_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt4_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt4_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt4_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt4_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt4_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt4_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt4_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt4_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt4_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt4_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt4_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt4_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt4_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt4_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt4_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt4_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt4_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt4_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt4_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt4_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt4_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt4_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt4_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt4_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt4_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt4_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt4_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt4_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt4_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt4_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt4_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt4_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt4_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt4_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt4_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt4_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt4_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt4_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt4_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[4] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt4_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[4] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt4_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt5_sd_pvld
  ) begin
    wt5_sd_pvld_w = wt_pre_sel[5] ? 1'b1 :
                    dat_pre_stripe_st[5] ? 1'b0 :
                    wt5_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt5_sd_pvld <= 1'b0;
  end else begin
  wt5_sd_pvld <= wt5_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5]) == 1'b1) begin
    wt5_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[5]) == 1'b0) begin
  end else begin
    wt5_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b1) begin
    wt5_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b0) begin
  end else begin
    wt5_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b1) begin
    wt5_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b0) begin
  end else begin
    wt5_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b1) begin
    wt5_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[5] & cfg_is_fp16_d1[71]) == 1'b0) begin
  end else begin
    wt5_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt5_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt5_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt5_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt5_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt5_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt5_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt5_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt5_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt5_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt5_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt5_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt5_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt5_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt5_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt5_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt5_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt5_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt5_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt5_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt5_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt5_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt5_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt5_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt5_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt5_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt5_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt5_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt5_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt5_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt5_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt5_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt5_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt5_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt5_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt5_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt5_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt5_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt5_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt5_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt5_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt5_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt5_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt5_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt5_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt5_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt5_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt5_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt5_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt5_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt5_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt5_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt5_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt5_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt5_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt5_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt5_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt5_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt5_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt5_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt5_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt5_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt5_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt5_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt5_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt5_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt5_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt5_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt5_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt5_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt5_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt5_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt5_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt5_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt5_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt5_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt5_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt5_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt5_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt5_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt5_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt5_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt5_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt5_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt5_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt5_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt5_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt5_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt5_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt5_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt5_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt5_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt5_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt5_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt5_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt5_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt5_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt5_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt5_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt5_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt5_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt5_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt5_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt5_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt5_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt5_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt5_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt5_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt5_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt5_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt5_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt5_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt5_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt5_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt5_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt5_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt5_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt5_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt5_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt5_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt5_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt5_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt5_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt5_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt5_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt5_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt5_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt5_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt5_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt5_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt5_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt5_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt5_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt5_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt5_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt5_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt5_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt5_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt5_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt5_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt5_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt5_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt5_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt5_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt5_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt5_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt5_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt5_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt5_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt5_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt5_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt5_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt5_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt5_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt5_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt5_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt5_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt5_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt5_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt5_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt5_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt5_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt5_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt5_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt5_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt5_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt5_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt5_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt5_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt5_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt5_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt5_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt5_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt5_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt5_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt5_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt5_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt5_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt5_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt5_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt5_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt5_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt5_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt5_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt5_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt5_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt5_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt5_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt5_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt5_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt5_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt5_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt5_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt5_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt5_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt5_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt5_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt5_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt5_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt5_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt5_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt5_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt5_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt5_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt5_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt5_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt5_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt5_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt5_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt5_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt5_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt5_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt5_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt5_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt5_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt5_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt5_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt5_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt5_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt5_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt5_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt5_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt5_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt5_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt5_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt5_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt5_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt5_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt5_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt5_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt5_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt5_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt5_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt5_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt5_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt5_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt5_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt5_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt5_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt5_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt5_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt5_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt5_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt5_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt5_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt5_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt5_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt5_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt5_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt5_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt5_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt5_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt5_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt5_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt5_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[5] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt5_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[5] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt5_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt6_sd_pvld
  ) begin
    wt6_sd_pvld_w = wt_pre_sel[6] ? 1'b1 :
                    dat_pre_stripe_st[6] ? 1'b0 :
                    wt6_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt6_sd_pvld <= 1'b0;
  end else begin
  wt6_sd_pvld <= wt6_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6]) == 1'b1) begin
    wt6_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[6]) == 1'b0) begin
  end else begin
    wt6_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b1) begin
    wt6_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b0) begin
  end else begin
    wt6_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b1) begin
    wt6_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b0) begin
  end else begin
    wt6_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b1) begin
    wt6_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[6] & cfg_is_fp16_d1[72]) == 1'b0) begin
  end else begin
    wt6_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt6_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt6_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt6_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt6_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt6_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt6_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt6_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt6_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt6_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt6_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt6_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt6_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt6_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt6_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt6_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt6_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt6_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt6_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt6_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt6_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt6_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt6_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt6_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt6_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt6_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt6_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt6_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt6_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt6_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt6_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt6_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt6_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt6_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt6_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt6_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt6_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt6_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt6_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt6_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt6_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt6_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt6_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt6_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt6_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt6_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt6_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt6_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt6_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt6_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt6_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt6_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt6_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt6_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt6_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt6_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt6_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt6_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt6_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt6_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt6_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt6_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt6_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt6_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt6_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt6_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt6_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt6_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt6_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt6_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt6_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt6_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt6_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt6_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt6_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt6_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt6_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt6_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt6_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt6_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt6_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt6_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt6_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt6_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt6_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt6_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt6_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt6_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt6_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt6_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt6_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt6_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt6_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt6_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt6_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt6_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt6_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt6_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt6_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt6_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt6_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt6_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt6_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt6_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt6_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt6_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt6_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt6_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt6_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt6_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt6_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt6_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt6_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt6_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt6_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt6_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt6_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt6_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt6_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt6_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt6_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt6_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt6_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt6_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt6_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt6_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt6_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt6_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt6_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt6_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt6_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt6_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt6_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt6_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt6_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt6_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt6_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt6_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt6_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt6_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt6_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt6_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt6_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt6_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt6_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt6_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt6_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt6_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt6_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt6_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt6_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt6_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt6_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt6_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt6_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt6_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt6_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt6_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt6_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt6_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt6_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt6_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt6_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt6_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt6_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt6_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt6_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt6_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt6_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt6_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt6_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt6_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt6_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt6_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt6_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt6_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt6_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt6_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt6_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt6_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt6_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt6_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt6_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt6_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt6_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt6_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt6_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt6_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt6_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt6_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt6_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt6_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt6_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt6_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt6_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt6_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt6_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt6_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt6_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt6_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt6_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt6_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt6_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt6_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt6_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt6_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt6_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt6_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt6_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt6_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt6_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt6_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt6_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt6_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt6_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt6_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt6_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt6_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt6_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt6_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt6_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt6_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt6_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt6_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt6_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt6_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt6_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt6_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt6_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt6_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt6_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt6_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt6_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt6_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt6_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt6_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt6_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt6_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt6_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt6_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt6_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt6_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt6_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt6_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt6_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt6_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt6_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt6_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt6_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt6_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt6_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt6_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt6_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt6_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt6_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[6] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt6_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[6] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt6_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  wt_pre_sel
  or dat_pre_stripe_st
  or wt7_sd_pvld
  ) begin
    wt7_sd_pvld_w = wt_pre_sel[7] ? 1'b1 :
                    dat_pre_stripe_st[7] ? 1'b0 :
                    wt7_sd_pvld;
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt7_sd_pvld <= 1'b0;
  end else begin
  wt7_sd_pvld <= wt7_sd_pvld_w;
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7]) == 1'b1) begin
    wt7_sd_nz <= wt_pre_nz;
  // VCS coverage off
  end else if ((wt_pre_sel[7]) == 1'b0) begin
  end else begin
    wt7_sd_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b1) begin
    wt7_sd_mask <= wt_pre_mask;
  // VCS coverage off
  end else if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b0) begin
  end else begin
    wt7_sd_mask <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b1) begin
    wt7_sd_exp <= wt_pre_exp;
  // VCS coverage off
  end else if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b0) begin
  end else begin
    wt7_sd_exp <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b1) begin
    wt7_sd_nan <= wt_pre_nan;
  // VCS coverage off
  end else if ((wt_pre_sel[7] & cfg_is_fp16_d1[73]) == 1'b0) begin
  end else begin
    wt7_sd_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b1) begin
    wt7_sd_data[7:0] <= wt_pre_data[7:0];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[0] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt7_sd_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b1) begin
    wt7_sd_data[15:8] <= wt_pre_data[15:8];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[1] | wt_pre_nan[0])) == 1'b0) begin
  end else begin
    wt7_sd_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b1) begin
    wt7_sd_data[23:16] <= wt_pre_data[23:16];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[2] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt7_sd_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b1) begin
    wt7_sd_data[31:24] <= wt_pre_data[31:24];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[3] | wt_pre_nan[1])) == 1'b0) begin
  end else begin
    wt7_sd_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b1) begin
    wt7_sd_data[39:32] <= wt_pre_data[39:32];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[4] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt7_sd_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b1) begin
    wt7_sd_data[47:40] <= wt_pre_data[47:40];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[5] | wt_pre_nan[2])) == 1'b0) begin
  end else begin
    wt7_sd_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b1) begin
    wt7_sd_data[55:48] <= wt_pre_data[55:48];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[6] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt7_sd_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b1) begin
    wt7_sd_data[63:56] <= wt_pre_data[63:56];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[7] | wt_pre_nan[3])) == 1'b0) begin
  end else begin
    wt7_sd_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b1) begin
    wt7_sd_data[71:64] <= wt_pre_data[71:64];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[8] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt7_sd_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b1) begin
    wt7_sd_data[79:72] <= wt_pre_data[79:72];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[9] | wt_pre_nan[4])) == 1'b0) begin
  end else begin
    wt7_sd_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b1) begin
    wt7_sd_data[87:80] <= wt_pre_data[87:80];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[10] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt7_sd_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b1) begin
    wt7_sd_data[95:88] <= wt_pre_data[95:88];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[11] | wt_pre_nan[5])) == 1'b0) begin
  end else begin
    wt7_sd_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b1) begin
    wt7_sd_data[103:96] <= wt_pre_data[103:96];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[12] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt7_sd_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b1) begin
    wt7_sd_data[111:104] <= wt_pre_data[111:104];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[13] | wt_pre_nan[6])) == 1'b0) begin
  end else begin
    wt7_sd_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b1) begin
    wt7_sd_data[119:112] <= wt_pre_data[119:112];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[14] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt7_sd_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b1) begin
    wt7_sd_data[127:120] <= wt_pre_data[127:120];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[15] | wt_pre_nan[7])) == 1'b0) begin
  end else begin
    wt7_sd_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b1) begin
    wt7_sd_data[135:128] <= wt_pre_data[135:128];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[16] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt7_sd_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b1) begin
    wt7_sd_data[143:136] <= wt_pre_data[143:136];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[17] | wt_pre_nan[8])) == 1'b0) begin
  end else begin
    wt7_sd_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b1) begin
    wt7_sd_data[151:144] <= wt_pre_data[151:144];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[18] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt7_sd_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b1) begin
    wt7_sd_data[159:152] <= wt_pre_data[159:152];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[19] | wt_pre_nan[9])) == 1'b0) begin
  end else begin
    wt7_sd_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b1) begin
    wt7_sd_data[167:160] <= wt_pre_data[167:160];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[20] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt7_sd_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b1) begin
    wt7_sd_data[175:168] <= wt_pre_data[175:168];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[21] | wt_pre_nan[10])) == 1'b0) begin
  end else begin
    wt7_sd_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b1) begin
    wt7_sd_data[183:176] <= wt_pre_data[183:176];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[22] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt7_sd_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b1) begin
    wt7_sd_data[191:184] <= wt_pre_data[191:184];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[23] | wt_pre_nan[11])) == 1'b0) begin
  end else begin
    wt7_sd_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b1) begin
    wt7_sd_data[199:192] <= wt_pre_data[199:192];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[24] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt7_sd_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b1) begin
    wt7_sd_data[207:200] <= wt_pre_data[207:200];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[25] | wt_pre_nan[12])) == 1'b0) begin
  end else begin
    wt7_sd_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b1) begin
    wt7_sd_data[215:208] <= wt_pre_data[215:208];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[26] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt7_sd_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b1) begin
    wt7_sd_data[223:216] <= wt_pre_data[223:216];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[27] | wt_pre_nan[13])) == 1'b0) begin
  end else begin
    wt7_sd_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b1) begin
    wt7_sd_data[231:224] <= wt_pre_data[231:224];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[28] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt7_sd_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b1) begin
    wt7_sd_data[239:232] <= wt_pre_data[239:232];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[29] | wt_pre_nan[14])) == 1'b0) begin
  end else begin
    wt7_sd_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b1) begin
    wt7_sd_data[247:240] <= wt_pre_data[247:240];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[30] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt7_sd_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b1) begin
    wt7_sd_data[255:248] <= wt_pre_data[255:248];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[31] | wt_pre_nan[15])) == 1'b0) begin
  end else begin
    wt7_sd_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b1) begin
    wt7_sd_data[263:256] <= wt_pre_data[263:256];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[32] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt7_sd_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b1) begin
    wt7_sd_data[271:264] <= wt_pre_data[271:264];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[33] | wt_pre_nan[16])) == 1'b0) begin
  end else begin
    wt7_sd_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b1) begin
    wt7_sd_data[279:272] <= wt_pre_data[279:272];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[34] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt7_sd_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b1) begin
    wt7_sd_data[287:280] <= wt_pre_data[287:280];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[35] | wt_pre_nan[17])) == 1'b0) begin
  end else begin
    wt7_sd_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b1) begin
    wt7_sd_data[295:288] <= wt_pre_data[295:288];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[36] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt7_sd_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b1) begin
    wt7_sd_data[303:296] <= wt_pre_data[303:296];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[37] | wt_pre_nan[18])) == 1'b0) begin
  end else begin
    wt7_sd_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b1) begin
    wt7_sd_data[311:304] <= wt_pre_data[311:304];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[38] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt7_sd_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b1) begin
    wt7_sd_data[319:312] <= wt_pre_data[319:312];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[39] | wt_pre_nan[19])) == 1'b0) begin
  end else begin
    wt7_sd_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b1) begin
    wt7_sd_data[327:320] <= wt_pre_data[327:320];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[40] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt7_sd_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b1) begin
    wt7_sd_data[335:328] <= wt_pre_data[335:328];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[41] | wt_pre_nan[20])) == 1'b0) begin
  end else begin
    wt7_sd_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b1) begin
    wt7_sd_data[343:336] <= wt_pre_data[343:336];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[42] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt7_sd_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b1) begin
    wt7_sd_data[351:344] <= wt_pre_data[351:344];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[43] | wt_pre_nan[21])) == 1'b0) begin
  end else begin
    wt7_sd_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b1) begin
    wt7_sd_data[359:352] <= wt_pre_data[359:352];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[44] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt7_sd_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b1) begin
    wt7_sd_data[367:360] <= wt_pre_data[367:360];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[45] | wt_pre_nan[22])) == 1'b0) begin
  end else begin
    wt7_sd_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b1) begin
    wt7_sd_data[375:368] <= wt_pre_data[375:368];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[46] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt7_sd_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b1) begin
    wt7_sd_data[383:376] <= wt_pre_data[383:376];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[47] | wt_pre_nan[23])) == 1'b0) begin
  end else begin
    wt7_sd_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b1) begin
    wt7_sd_data[391:384] <= wt_pre_data[391:384];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[48] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt7_sd_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b1) begin
    wt7_sd_data[399:392] <= wt_pre_data[399:392];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[49] | wt_pre_nan[24])) == 1'b0) begin
  end else begin
    wt7_sd_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b1) begin
    wt7_sd_data[407:400] <= wt_pre_data[407:400];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[50] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt7_sd_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b1) begin
    wt7_sd_data[415:408] <= wt_pre_data[415:408];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[51] | wt_pre_nan[25])) == 1'b0) begin
  end else begin
    wt7_sd_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b1) begin
    wt7_sd_data[423:416] <= wt_pre_data[423:416];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[52] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt7_sd_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b1) begin
    wt7_sd_data[431:424] <= wt_pre_data[431:424];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[53] | wt_pre_nan[26])) == 1'b0) begin
  end else begin
    wt7_sd_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b1) begin
    wt7_sd_data[439:432] <= wt_pre_data[439:432];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[54] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt7_sd_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b1) begin
    wt7_sd_data[447:440] <= wt_pre_data[447:440];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[55] | wt_pre_nan[27])) == 1'b0) begin
  end else begin
    wt7_sd_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b1) begin
    wt7_sd_data[455:448] <= wt_pre_data[455:448];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[56] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt7_sd_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b1) begin
    wt7_sd_data[463:456] <= wt_pre_data[463:456];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[57] | wt_pre_nan[28])) == 1'b0) begin
  end else begin
    wt7_sd_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b1) begin
    wt7_sd_data[471:464] <= wt_pre_data[471:464];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[58] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt7_sd_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b1) begin
    wt7_sd_data[479:472] <= wt_pre_data[479:472];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[59] | wt_pre_nan[29])) == 1'b0) begin
  end else begin
    wt7_sd_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b1) begin
    wt7_sd_data[487:480] <= wt_pre_data[487:480];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[60] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt7_sd_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b1) begin
    wt7_sd_data[495:488] <= wt_pre_data[495:488];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[61] | wt_pre_nan[30])) == 1'b0) begin
  end else begin
    wt7_sd_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b1) begin
    wt7_sd_data[503:496] <= wt_pre_data[503:496];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[62] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt7_sd_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b1) begin
    wt7_sd_data[511:504] <= wt_pre_data[511:504];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[63] | wt_pre_nan[31])) == 1'b0) begin
  end else begin
    wt7_sd_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b1) begin
    wt7_sd_data[519:512] <= wt_pre_data[519:512];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[64] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt7_sd_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b1) begin
    wt7_sd_data[527:520] <= wt_pre_data[527:520];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[65] | wt_pre_nan[32])) == 1'b0) begin
  end else begin
    wt7_sd_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b1) begin
    wt7_sd_data[535:528] <= wt_pre_data[535:528];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[66] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt7_sd_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b1) begin
    wt7_sd_data[543:536] <= wt_pre_data[543:536];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[67] | wt_pre_nan[33])) == 1'b0) begin
  end else begin
    wt7_sd_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b1) begin
    wt7_sd_data[551:544] <= wt_pre_data[551:544];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[68] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt7_sd_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b1) begin
    wt7_sd_data[559:552] <= wt_pre_data[559:552];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[69] | wt_pre_nan[34])) == 1'b0) begin
  end else begin
    wt7_sd_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b1) begin
    wt7_sd_data[567:560] <= wt_pre_data[567:560];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[70] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt7_sd_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b1) begin
    wt7_sd_data[575:568] <= wt_pre_data[575:568];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[71] | wt_pre_nan[35])) == 1'b0) begin
  end else begin
    wt7_sd_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b1) begin
    wt7_sd_data[583:576] <= wt_pre_data[583:576];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[72] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt7_sd_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b1) begin
    wt7_sd_data[591:584] <= wt_pre_data[591:584];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[73] | wt_pre_nan[36])) == 1'b0) begin
  end else begin
    wt7_sd_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b1) begin
    wt7_sd_data[599:592] <= wt_pre_data[599:592];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[74] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt7_sd_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b1) begin
    wt7_sd_data[607:600] <= wt_pre_data[607:600];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[75] | wt_pre_nan[37])) == 1'b0) begin
  end else begin
    wt7_sd_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b1) begin
    wt7_sd_data[615:608] <= wt_pre_data[615:608];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[76] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt7_sd_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b1) begin
    wt7_sd_data[623:616] <= wt_pre_data[623:616];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[77] | wt_pre_nan[38])) == 1'b0) begin
  end else begin
    wt7_sd_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b1) begin
    wt7_sd_data[631:624] <= wt_pre_data[631:624];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[78] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt7_sd_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b1) begin
    wt7_sd_data[639:632] <= wt_pre_data[639:632];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[79] | wt_pre_nan[39])) == 1'b0) begin
  end else begin
    wt7_sd_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b1) begin
    wt7_sd_data[647:640] <= wt_pre_data[647:640];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[80] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt7_sd_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b1) begin
    wt7_sd_data[655:648] <= wt_pre_data[655:648];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[81] | wt_pre_nan[40])) == 1'b0) begin
  end else begin
    wt7_sd_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b1) begin
    wt7_sd_data[663:656] <= wt_pre_data[663:656];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[82] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt7_sd_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b1) begin
    wt7_sd_data[671:664] <= wt_pre_data[671:664];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[83] | wt_pre_nan[41])) == 1'b0) begin
  end else begin
    wt7_sd_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b1) begin
    wt7_sd_data[679:672] <= wt_pre_data[679:672];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[84] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt7_sd_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b1) begin
    wt7_sd_data[687:680] <= wt_pre_data[687:680];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[85] | wt_pre_nan[42])) == 1'b0) begin
  end else begin
    wt7_sd_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b1) begin
    wt7_sd_data[695:688] <= wt_pre_data[695:688];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[86] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt7_sd_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b1) begin
    wt7_sd_data[703:696] <= wt_pre_data[703:696];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[87] | wt_pre_nan[43])) == 1'b0) begin
  end else begin
    wt7_sd_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b1) begin
    wt7_sd_data[711:704] <= wt_pre_data[711:704];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[88] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt7_sd_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b1) begin
    wt7_sd_data[719:712] <= wt_pre_data[719:712];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[89] | wt_pre_nan[44])) == 1'b0) begin
  end else begin
    wt7_sd_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b1) begin
    wt7_sd_data[727:720] <= wt_pre_data[727:720];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[90] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt7_sd_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b1) begin
    wt7_sd_data[735:728] <= wt_pre_data[735:728];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[91] | wt_pre_nan[45])) == 1'b0) begin
  end else begin
    wt7_sd_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b1) begin
    wt7_sd_data[743:736] <= wt_pre_data[743:736];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[92] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt7_sd_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b1) begin
    wt7_sd_data[751:744] <= wt_pre_data[751:744];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[93] | wt_pre_nan[46])) == 1'b0) begin
  end else begin
    wt7_sd_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b1) begin
    wt7_sd_data[759:752] <= wt_pre_data[759:752];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[94] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt7_sd_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b1) begin
    wt7_sd_data[767:760] <= wt_pre_data[767:760];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[95] | wt_pre_nan[47])) == 1'b0) begin
  end else begin
    wt7_sd_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b1) begin
    wt7_sd_data[775:768] <= wt_pre_data[775:768];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[96] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt7_sd_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b1) begin
    wt7_sd_data[783:776] <= wt_pre_data[783:776];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[97] | wt_pre_nan[48])) == 1'b0) begin
  end else begin
    wt7_sd_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b1) begin
    wt7_sd_data[791:784] <= wt_pre_data[791:784];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[98] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt7_sd_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b1) begin
    wt7_sd_data[799:792] <= wt_pre_data[799:792];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[99] | wt_pre_nan[49])) == 1'b0) begin
  end else begin
    wt7_sd_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b1) begin
    wt7_sd_data[807:800] <= wt_pre_data[807:800];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[100] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt7_sd_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b1) begin
    wt7_sd_data[815:808] <= wt_pre_data[815:808];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[101] | wt_pre_nan[50])) == 1'b0) begin
  end else begin
    wt7_sd_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b1) begin
    wt7_sd_data[823:816] <= wt_pre_data[823:816];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[102] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt7_sd_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b1) begin
    wt7_sd_data[831:824] <= wt_pre_data[831:824];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[103] | wt_pre_nan[51])) == 1'b0) begin
  end else begin
    wt7_sd_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b1) begin
    wt7_sd_data[839:832] <= wt_pre_data[839:832];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[104] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt7_sd_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b1) begin
    wt7_sd_data[847:840] <= wt_pre_data[847:840];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[105] | wt_pre_nan[52])) == 1'b0) begin
  end else begin
    wt7_sd_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b1) begin
    wt7_sd_data[855:848] <= wt_pre_data[855:848];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[106] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt7_sd_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b1) begin
    wt7_sd_data[863:856] <= wt_pre_data[863:856];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[107] | wt_pre_nan[53])) == 1'b0) begin
  end else begin
    wt7_sd_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b1) begin
    wt7_sd_data[871:864] <= wt_pre_data[871:864];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[108] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt7_sd_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b1) begin
    wt7_sd_data[879:872] <= wt_pre_data[879:872];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[109] | wt_pre_nan[54])) == 1'b0) begin
  end else begin
    wt7_sd_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b1) begin
    wt7_sd_data[887:880] <= wt_pre_data[887:880];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[110] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt7_sd_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b1) begin
    wt7_sd_data[895:888] <= wt_pre_data[895:888];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[111] | wt_pre_nan[55])) == 1'b0) begin
  end else begin
    wt7_sd_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b1) begin
    wt7_sd_data[903:896] <= wt_pre_data[903:896];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[112] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt7_sd_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b1) begin
    wt7_sd_data[911:904] <= wt_pre_data[911:904];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[113] | wt_pre_nan[56])) == 1'b0) begin
  end else begin
    wt7_sd_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b1) begin
    wt7_sd_data[919:912] <= wt_pre_data[919:912];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[114] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt7_sd_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b1) begin
    wt7_sd_data[927:920] <= wt_pre_data[927:920];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[115] | wt_pre_nan[57])) == 1'b0) begin
  end else begin
    wt7_sd_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b1) begin
    wt7_sd_data[935:928] <= wt_pre_data[935:928];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[116] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt7_sd_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b1) begin
    wt7_sd_data[943:936] <= wt_pre_data[943:936];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[117] | wt_pre_nan[58])) == 1'b0) begin
  end else begin
    wt7_sd_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b1) begin
    wt7_sd_data[951:944] <= wt_pre_data[951:944];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[118] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt7_sd_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b1) begin
    wt7_sd_data[959:952] <= wt_pre_data[959:952];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[119] | wt_pre_nan[59])) == 1'b0) begin
  end else begin
    wt7_sd_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b1) begin
    wt7_sd_data[967:960] <= wt_pre_data[967:960];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[120] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt7_sd_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b1) begin
    wt7_sd_data[975:968] <= wt_pre_data[975:968];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[121] | wt_pre_nan[60])) == 1'b0) begin
  end else begin
    wt7_sd_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b1) begin
    wt7_sd_data[983:976] <= wt_pre_data[983:976];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[122] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt7_sd_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b1) begin
    wt7_sd_data[991:984] <= wt_pre_data[991:984];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[123] | wt_pre_nan[61])) == 1'b0) begin
  end else begin
    wt7_sd_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b1) begin
    wt7_sd_data[999:992] <= wt_pre_data[999:992];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[124] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt7_sd_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b1) begin
    wt7_sd_data[1007:1000] <= wt_pre_data[1007:1000];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[125] | wt_pre_nan[62])) == 1'b0) begin
  end else begin
    wt7_sd_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b1) begin
    wt7_sd_data[1015:1008] <= wt_pre_data[1015:1008];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[126] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt7_sd_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((wt_pre_sel[7] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b1) begin
    wt7_sd_data[1023:1016] <= wt_pre_data[1023:1016];
  // VCS coverage off
  end else if ((wt_pre_sel[7] & (wt_pre_nz[127] | wt_pre_nan[63])) == 1'b0) begin
  end else begin
    wt7_sd_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end










always @(
  dat_pre_stripe_st
  or wt0_sd_pvld
  or dat_actv_stripe_end
  or wt0_actv_vld
  ) begin
    wt0_actv_pvld_w = dat_pre_stripe_st[0] ? wt0_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt0_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt0_actv_vld <= 1'b0;
  end else begin
  wt0_actv_vld <= wt0_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt0_actv_pvld <= {104{1'b0}};
  end else begin
  wt0_actv_pvld <= {104{wt0_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_nz <= wt0_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w & cfg_is_fp16_d1[74]) == 1'b1) begin
    wt0_actv_nan <= wt0_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w & cfg_is_fp16_d1[74]) == 1'b0) begin
  end else begin
    wt0_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[7:0] <= {8{(wt0_sd_nz[0] | wt0_sd_nan[0])}} & wt0_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[15:8] <= {8{(wt0_sd_nz[1] | wt0_sd_nan[0])}} & wt0_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[23:16] <= {8{(wt0_sd_nz[2] | wt0_sd_nan[1])}} & wt0_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[31:24] <= {8{(wt0_sd_nz[3] | wt0_sd_nan[1])}} & wt0_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[39:32] <= {8{(wt0_sd_nz[4] | wt0_sd_nan[2])}} & wt0_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[47:40] <= {8{(wt0_sd_nz[5] | wt0_sd_nan[2])}} & wt0_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[55:48] <= {8{(wt0_sd_nz[6] | wt0_sd_nan[3])}} & wt0_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[63:56] <= {8{(wt0_sd_nz[7] | wt0_sd_nan[3])}} & wt0_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[71:64] <= {8{(wt0_sd_nz[8] | wt0_sd_nan[4])}} & wt0_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[79:72] <= {8{(wt0_sd_nz[9] | wt0_sd_nan[4])}} & wt0_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[87:80] <= {8{(wt0_sd_nz[10] | wt0_sd_nan[5])}} & wt0_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[95:88] <= {8{(wt0_sd_nz[11] | wt0_sd_nan[5])}} & wt0_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[103:96] <= {8{(wt0_sd_nz[12] | wt0_sd_nan[6])}} & wt0_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[111:104] <= {8{(wt0_sd_nz[13] | wt0_sd_nan[6])}} & wt0_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[119:112] <= {8{(wt0_sd_nz[14] | wt0_sd_nan[7])}} & wt0_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[127:120] <= {8{(wt0_sd_nz[15] | wt0_sd_nan[7])}} & wt0_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[135:128] <= {8{(wt0_sd_nz[16] | wt0_sd_nan[8])}} & wt0_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[143:136] <= {8{(wt0_sd_nz[17] | wt0_sd_nan[8])}} & wt0_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[151:144] <= {8{(wt0_sd_nz[18] | wt0_sd_nan[9])}} & wt0_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[159:152] <= {8{(wt0_sd_nz[19] | wt0_sd_nan[9])}} & wt0_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[167:160] <= {8{(wt0_sd_nz[20] | wt0_sd_nan[10])}} & wt0_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[175:168] <= {8{(wt0_sd_nz[21] | wt0_sd_nan[10])}} & wt0_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[183:176] <= {8{(wt0_sd_nz[22] | wt0_sd_nan[11])}} & wt0_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[191:184] <= {8{(wt0_sd_nz[23] | wt0_sd_nan[11])}} & wt0_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[199:192] <= {8{(wt0_sd_nz[24] | wt0_sd_nan[12])}} & wt0_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[207:200] <= {8{(wt0_sd_nz[25] | wt0_sd_nan[12])}} & wt0_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[215:208] <= {8{(wt0_sd_nz[26] | wt0_sd_nan[13])}} & wt0_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[223:216] <= {8{(wt0_sd_nz[27] | wt0_sd_nan[13])}} & wt0_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[231:224] <= {8{(wt0_sd_nz[28] | wt0_sd_nan[14])}} & wt0_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[239:232] <= {8{(wt0_sd_nz[29] | wt0_sd_nan[14])}} & wt0_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[247:240] <= {8{(wt0_sd_nz[30] | wt0_sd_nan[15])}} & wt0_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[255:248] <= {8{(wt0_sd_nz[31] | wt0_sd_nan[15])}} & wt0_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[263:256] <= {8{(wt0_sd_nz[32] | wt0_sd_nan[16])}} & wt0_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[271:264] <= {8{(wt0_sd_nz[33] | wt0_sd_nan[16])}} & wt0_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[279:272] <= {8{(wt0_sd_nz[34] | wt0_sd_nan[17])}} & wt0_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[287:280] <= {8{(wt0_sd_nz[35] | wt0_sd_nan[17])}} & wt0_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[295:288] <= {8{(wt0_sd_nz[36] | wt0_sd_nan[18])}} & wt0_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[303:296] <= {8{(wt0_sd_nz[37] | wt0_sd_nan[18])}} & wt0_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[311:304] <= {8{(wt0_sd_nz[38] | wt0_sd_nan[19])}} & wt0_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[319:312] <= {8{(wt0_sd_nz[39] | wt0_sd_nan[19])}} & wt0_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[327:320] <= {8{(wt0_sd_nz[40] | wt0_sd_nan[20])}} & wt0_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[335:328] <= {8{(wt0_sd_nz[41] | wt0_sd_nan[20])}} & wt0_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[343:336] <= {8{(wt0_sd_nz[42] | wt0_sd_nan[21])}} & wt0_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[351:344] <= {8{(wt0_sd_nz[43] | wt0_sd_nan[21])}} & wt0_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[359:352] <= {8{(wt0_sd_nz[44] | wt0_sd_nan[22])}} & wt0_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[367:360] <= {8{(wt0_sd_nz[45] | wt0_sd_nan[22])}} & wt0_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[375:368] <= {8{(wt0_sd_nz[46] | wt0_sd_nan[23])}} & wt0_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[383:376] <= {8{(wt0_sd_nz[47] | wt0_sd_nan[23])}} & wt0_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[391:384] <= {8{(wt0_sd_nz[48] | wt0_sd_nan[24])}} & wt0_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[399:392] <= {8{(wt0_sd_nz[49] | wt0_sd_nan[24])}} & wt0_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[407:400] <= {8{(wt0_sd_nz[50] | wt0_sd_nan[25])}} & wt0_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[415:408] <= {8{(wt0_sd_nz[51] | wt0_sd_nan[25])}} & wt0_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[423:416] <= {8{(wt0_sd_nz[52] | wt0_sd_nan[26])}} & wt0_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[431:424] <= {8{(wt0_sd_nz[53] | wt0_sd_nan[26])}} & wt0_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[439:432] <= {8{(wt0_sd_nz[54] | wt0_sd_nan[27])}} & wt0_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[447:440] <= {8{(wt0_sd_nz[55] | wt0_sd_nan[27])}} & wt0_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[455:448] <= {8{(wt0_sd_nz[56] | wt0_sd_nan[28])}} & wt0_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[463:456] <= {8{(wt0_sd_nz[57] | wt0_sd_nan[28])}} & wt0_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[471:464] <= {8{(wt0_sd_nz[58] | wt0_sd_nan[29])}} & wt0_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[479:472] <= {8{(wt0_sd_nz[59] | wt0_sd_nan[29])}} & wt0_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[487:480] <= {8{(wt0_sd_nz[60] | wt0_sd_nan[30])}} & wt0_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[495:488] <= {8{(wt0_sd_nz[61] | wt0_sd_nan[30])}} & wt0_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[503:496] <= {8{(wt0_sd_nz[62] | wt0_sd_nan[31])}} & wt0_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[511:504] <= {8{(wt0_sd_nz[63] | wt0_sd_nan[31])}} & wt0_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[519:512] <= {8{(wt0_sd_nz[64] | wt0_sd_nan[32])}} & wt0_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[527:520] <= {8{(wt0_sd_nz[65] | wt0_sd_nan[32])}} & wt0_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[535:528] <= {8{(wt0_sd_nz[66] | wt0_sd_nan[33])}} & wt0_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[543:536] <= {8{(wt0_sd_nz[67] | wt0_sd_nan[33])}} & wt0_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[551:544] <= {8{(wt0_sd_nz[68] | wt0_sd_nan[34])}} & wt0_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[559:552] <= {8{(wt0_sd_nz[69] | wt0_sd_nan[34])}} & wt0_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[567:560] <= {8{(wt0_sd_nz[70] | wt0_sd_nan[35])}} & wt0_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[575:568] <= {8{(wt0_sd_nz[71] | wt0_sd_nan[35])}} & wt0_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[583:576] <= {8{(wt0_sd_nz[72] | wt0_sd_nan[36])}} & wt0_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[591:584] <= {8{(wt0_sd_nz[73] | wt0_sd_nan[36])}} & wt0_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[599:592] <= {8{(wt0_sd_nz[74] | wt0_sd_nan[37])}} & wt0_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[607:600] <= {8{(wt0_sd_nz[75] | wt0_sd_nan[37])}} & wt0_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[615:608] <= {8{(wt0_sd_nz[76] | wt0_sd_nan[38])}} & wt0_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[623:616] <= {8{(wt0_sd_nz[77] | wt0_sd_nan[38])}} & wt0_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[631:624] <= {8{(wt0_sd_nz[78] | wt0_sd_nan[39])}} & wt0_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[639:632] <= {8{(wt0_sd_nz[79] | wt0_sd_nan[39])}} & wt0_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[647:640] <= {8{(wt0_sd_nz[80] | wt0_sd_nan[40])}} & wt0_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[655:648] <= {8{(wt0_sd_nz[81] | wt0_sd_nan[40])}} & wt0_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[663:656] <= {8{(wt0_sd_nz[82] | wt0_sd_nan[41])}} & wt0_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[671:664] <= {8{(wt0_sd_nz[83] | wt0_sd_nan[41])}} & wt0_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[679:672] <= {8{(wt0_sd_nz[84] | wt0_sd_nan[42])}} & wt0_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[687:680] <= {8{(wt0_sd_nz[85] | wt0_sd_nan[42])}} & wt0_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[695:688] <= {8{(wt0_sd_nz[86] | wt0_sd_nan[43])}} & wt0_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[703:696] <= {8{(wt0_sd_nz[87] | wt0_sd_nan[43])}} & wt0_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[711:704] <= {8{(wt0_sd_nz[88] | wt0_sd_nan[44])}} & wt0_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[719:712] <= {8{(wt0_sd_nz[89] | wt0_sd_nan[44])}} & wt0_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[727:720] <= {8{(wt0_sd_nz[90] | wt0_sd_nan[45])}} & wt0_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[735:728] <= {8{(wt0_sd_nz[91] | wt0_sd_nan[45])}} & wt0_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[743:736] <= {8{(wt0_sd_nz[92] | wt0_sd_nan[46])}} & wt0_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[751:744] <= {8{(wt0_sd_nz[93] | wt0_sd_nan[46])}} & wt0_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[759:752] <= {8{(wt0_sd_nz[94] | wt0_sd_nan[47])}} & wt0_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[767:760] <= {8{(wt0_sd_nz[95] | wt0_sd_nan[47])}} & wt0_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[775:768] <= {8{(wt0_sd_nz[96] | wt0_sd_nan[48])}} & wt0_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[783:776] <= {8{(wt0_sd_nz[97] | wt0_sd_nan[48])}} & wt0_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[791:784] <= {8{(wt0_sd_nz[98] | wt0_sd_nan[49])}} & wt0_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[799:792] <= {8{(wt0_sd_nz[99] | wt0_sd_nan[49])}} & wt0_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[807:800] <= {8{(wt0_sd_nz[100] | wt0_sd_nan[50])}} & wt0_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[815:808] <= {8{(wt0_sd_nz[101] | wt0_sd_nan[50])}} & wt0_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[823:816] <= {8{(wt0_sd_nz[102] | wt0_sd_nan[51])}} & wt0_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[831:824] <= {8{(wt0_sd_nz[103] | wt0_sd_nan[51])}} & wt0_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[839:832] <= {8{(wt0_sd_nz[104] | wt0_sd_nan[52])}} & wt0_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[847:840] <= {8{(wt0_sd_nz[105] | wt0_sd_nan[52])}} & wt0_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[855:848] <= {8{(wt0_sd_nz[106] | wt0_sd_nan[53])}} & wt0_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[863:856] <= {8{(wt0_sd_nz[107] | wt0_sd_nan[53])}} & wt0_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[871:864] <= {8{(wt0_sd_nz[108] | wt0_sd_nan[54])}} & wt0_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[879:872] <= {8{(wt0_sd_nz[109] | wt0_sd_nan[54])}} & wt0_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[887:880] <= {8{(wt0_sd_nz[110] | wt0_sd_nan[55])}} & wt0_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[895:888] <= {8{(wt0_sd_nz[111] | wt0_sd_nan[55])}} & wt0_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[903:896] <= {8{(wt0_sd_nz[112] | wt0_sd_nan[56])}} & wt0_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[911:904] <= {8{(wt0_sd_nz[113] | wt0_sd_nan[56])}} & wt0_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[919:912] <= {8{(wt0_sd_nz[114] | wt0_sd_nan[57])}} & wt0_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[927:920] <= {8{(wt0_sd_nz[115] | wt0_sd_nan[57])}} & wt0_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[935:928] <= {8{(wt0_sd_nz[116] | wt0_sd_nan[58])}} & wt0_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[943:936] <= {8{(wt0_sd_nz[117] | wt0_sd_nan[58])}} & wt0_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[951:944] <= {8{(wt0_sd_nz[118] | wt0_sd_nan[59])}} & wt0_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[959:952] <= {8{(wt0_sd_nz[119] | wt0_sd_nan[59])}} & wt0_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[967:960] <= {8{(wt0_sd_nz[120] | wt0_sd_nan[60])}} & wt0_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[975:968] <= {8{(wt0_sd_nz[121] | wt0_sd_nan[60])}} & wt0_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[983:976] <= {8{(wt0_sd_nz[122] | wt0_sd_nan[61])}} & wt0_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[991:984] <= {8{(wt0_sd_nz[123] | wt0_sd_nan[61])}} & wt0_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[999:992] <= {8{(wt0_sd_nz[124] | wt0_sd_nan[62])}} & wt0_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[1007:1000] <= {8{(wt0_sd_nz[125] | wt0_sd_nan[62])}} & wt0_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[1015:1008] <= {8{(wt0_sd_nz[126] | wt0_sd_nan[63])}} & wt0_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b1) begin
    wt0_actv_data[1023:1016] <= {8{(wt0_sd_nz[127] | wt0_sd_nan[63])}} & wt0_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[0] & wt0_actv_pvld_w) == 1'b0) begin
  end else begin
    wt0_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt1_sd_pvld
  or dat_actv_stripe_end
  or wt1_actv_vld
  ) begin
    wt1_actv_pvld_w = dat_pre_stripe_st[1] ? wt1_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt1_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt1_actv_vld <= 1'b0;
  end else begin
  wt1_actv_vld <= wt1_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt1_actv_pvld <= {104{1'b0}};
  end else begin
  wt1_actv_pvld <= {104{wt1_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_nz <= wt1_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w & cfg_is_fp16_d1[75]) == 1'b1) begin
    wt1_actv_nan <= wt1_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w & cfg_is_fp16_d1[75]) == 1'b0) begin
  end else begin
    wt1_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[7:0] <= {8{(wt1_sd_nz[0] | wt1_sd_nan[0])}} & wt1_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[15:8] <= {8{(wt1_sd_nz[1] | wt1_sd_nan[0])}} & wt1_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[23:16] <= {8{(wt1_sd_nz[2] | wt1_sd_nan[1])}} & wt1_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[31:24] <= {8{(wt1_sd_nz[3] | wt1_sd_nan[1])}} & wt1_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[39:32] <= {8{(wt1_sd_nz[4] | wt1_sd_nan[2])}} & wt1_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[47:40] <= {8{(wt1_sd_nz[5] | wt1_sd_nan[2])}} & wt1_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[55:48] <= {8{(wt1_sd_nz[6] | wt1_sd_nan[3])}} & wt1_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[63:56] <= {8{(wt1_sd_nz[7] | wt1_sd_nan[3])}} & wt1_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[71:64] <= {8{(wt1_sd_nz[8] | wt1_sd_nan[4])}} & wt1_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[79:72] <= {8{(wt1_sd_nz[9] | wt1_sd_nan[4])}} & wt1_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[87:80] <= {8{(wt1_sd_nz[10] | wt1_sd_nan[5])}} & wt1_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[95:88] <= {8{(wt1_sd_nz[11] | wt1_sd_nan[5])}} & wt1_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[103:96] <= {8{(wt1_sd_nz[12] | wt1_sd_nan[6])}} & wt1_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[111:104] <= {8{(wt1_sd_nz[13] | wt1_sd_nan[6])}} & wt1_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[119:112] <= {8{(wt1_sd_nz[14] | wt1_sd_nan[7])}} & wt1_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[127:120] <= {8{(wt1_sd_nz[15] | wt1_sd_nan[7])}} & wt1_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[135:128] <= {8{(wt1_sd_nz[16] | wt1_sd_nan[8])}} & wt1_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[143:136] <= {8{(wt1_sd_nz[17] | wt1_sd_nan[8])}} & wt1_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[151:144] <= {8{(wt1_sd_nz[18] | wt1_sd_nan[9])}} & wt1_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[159:152] <= {8{(wt1_sd_nz[19] | wt1_sd_nan[9])}} & wt1_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[167:160] <= {8{(wt1_sd_nz[20] | wt1_sd_nan[10])}} & wt1_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[175:168] <= {8{(wt1_sd_nz[21] | wt1_sd_nan[10])}} & wt1_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[183:176] <= {8{(wt1_sd_nz[22] | wt1_sd_nan[11])}} & wt1_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[191:184] <= {8{(wt1_sd_nz[23] | wt1_sd_nan[11])}} & wt1_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[199:192] <= {8{(wt1_sd_nz[24] | wt1_sd_nan[12])}} & wt1_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[207:200] <= {8{(wt1_sd_nz[25] | wt1_sd_nan[12])}} & wt1_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[215:208] <= {8{(wt1_sd_nz[26] | wt1_sd_nan[13])}} & wt1_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[223:216] <= {8{(wt1_sd_nz[27] | wt1_sd_nan[13])}} & wt1_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[231:224] <= {8{(wt1_sd_nz[28] | wt1_sd_nan[14])}} & wt1_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[239:232] <= {8{(wt1_sd_nz[29] | wt1_sd_nan[14])}} & wt1_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[247:240] <= {8{(wt1_sd_nz[30] | wt1_sd_nan[15])}} & wt1_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[255:248] <= {8{(wt1_sd_nz[31] | wt1_sd_nan[15])}} & wt1_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[263:256] <= {8{(wt1_sd_nz[32] | wt1_sd_nan[16])}} & wt1_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[271:264] <= {8{(wt1_sd_nz[33] | wt1_sd_nan[16])}} & wt1_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[279:272] <= {8{(wt1_sd_nz[34] | wt1_sd_nan[17])}} & wt1_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[287:280] <= {8{(wt1_sd_nz[35] | wt1_sd_nan[17])}} & wt1_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[295:288] <= {8{(wt1_sd_nz[36] | wt1_sd_nan[18])}} & wt1_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[303:296] <= {8{(wt1_sd_nz[37] | wt1_sd_nan[18])}} & wt1_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[311:304] <= {8{(wt1_sd_nz[38] | wt1_sd_nan[19])}} & wt1_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[319:312] <= {8{(wt1_sd_nz[39] | wt1_sd_nan[19])}} & wt1_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[327:320] <= {8{(wt1_sd_nz[40] | wt1_sd_nan[20])}} & wt1_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[335:328] <= {8{(wt1_sd_nz[41] | wt1_sd_nan[20])}} & wt1_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[343:336] <= {8{(wt1_sd_nz[42] | wt1_sd_nan[21])}} & wt1_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[351:344] <= {8{(wt1_sd_nz[43] | wt1_sd_nan[21])}} & wt1_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[359:352] <= {8{(wt1_sd_nz[44] | wt1_sd_nan[22])}} & wt1_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[367:360] <= {8{(wt1_sd_nz[45] | wt1_sd_nan[22])}} & wt1_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[375:368] <= {8{(wt1_sd_nz[46] | wt1_sd_nan[23])}} & wt1_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[383:376] <= {8{(wt1_sd_nz[47] | wt1_sd_nan[23])}} & wt1_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[391:384] <= {8{(wt1_sd_nz[48] | wt1_sd_nan[24])}} & wt1_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[399:392] <= {8{(wt1_sd_nz[49] | wt1_sd_nan[24])}} & wt1_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[407:400] <= {8{(wt1_sd_nz[50] | wt1_sd_nan[25])}} & wt1_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[415:408] <= {8{(wt1_sd_nz[51] | wt1_sd_nan[25])}} & wt1_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[423:416] <= {8{(wt1_sd_nz[52] | wt1_sd_nan[26])}} & wt1_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[431:424] <= {8{(wt1_sd_nz[53] | wt1_sd_nan[26])}} & wt1_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[439:432] <= {8{(wt1_sd_nz[54] | wt1_sd_nan[27])}} & wt1_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[447:440] <= {8{(wt1_sd_nz[55] | wt1_sd_nan[27])}} & wt1_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[455:448] <= {8{(wt1_sd_nz[56] | wt1_sd_nan[28])}} & wt1_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[463:456] <= {8{(wt1_sd_nz[57] | wt1_sd_nan[28])}} & wt1_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[471:464] <= {8{(wt1_sd_nz[58] | wt1_sd_nan[29])}} & wt1_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[479:472] <= {8{(wt1_sd_nz[59] | wt1_sd_nan[29])}} & wt1_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[487:480] <= {8{(wt1_sd_nz[60] | wt1_sd_nan[30])}} & wt1_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[495:488] <= {8{(wt1_sd_nz[61] | wt1_sd_nan[30])}} & wt1_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[503:496] <= {8{(wt1_sd_nz[62] | wt1_sd_nan[31])}} & wt1_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[511:504] <= {8{(wt1_sd_nz[63] | wt1_sd_nan[31])}} & wt1_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[519:512] <= {8{(wt1_sd_nz[64] | wt1_sd_nan[32])}} & wt1_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[527:520] <= {8{(wt1_sd_nz[65] | wt1_sd_nan[32])}} & wt1_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[535:528] <= {8{(wt1_sd_nz[66] | wt1_sd_nan[33])}} & wt1_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[543:536] <= {8{(wt1_sd_nz[67] | wt1_sd_nan[33])}} & wt1_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[551:544] <= {8{(wt1_sd_nz[68] | wt1_sd_nan[34])}} & wt1_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[559:552] <= {8{(wt1_sd_nz[69] | wt1_sd_nan[34])}} & wt1_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[567:560] <= {8{(wt1_sd_nz[70] | wt1_sd_nan[35])}} & wt1_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[575:568] <= {8{(wt1_sd_nz[71] | wt1_sd_nan[35])}} & wt1_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[583:576] <= {8{(wt1_sd_nz[72] | wt1_sd_nan[36])}} & wt1_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[591:584] <= {8{(wt1_sd_nz[73] | wt1_sd_nan[36])}} & wt1_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[599:592] <= {8{(wt1_sd_nz[74] | wt1_sd_nan[37])}} & wt1_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[607:600] <= {8{(wt1_sd_nz[75] | wt1_sd_nan[37])}} & wt1_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[615:608] <= {8{(wt1_sd_nz[76] | wt1_sd_nan[38])}} & wt1_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[623:616] <= {8{(wt1_sd_nz[77] | wt1_sd_nan[38])}} & wt1_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[631:624] <= {8{(wt1_sd_nz[78] | wt1_sd_nan[39])}} & wt1_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[639:632] <= {8{(wt1_sd_nz[79] | wt1_sd_nan[39])}} & wt1_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[647:640] <= {8{(wt1_sd_nz[80] | wt1_sd_nan[40])}} & wt1_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[655:648] <= {8{(wt1_sd_nz[81] | wt1_sd_nan[40])}} & wt1_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[663:656] <= {8{(wt1_sd_nz[82] | wt1_sd_nan[41])}} & wt1_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[671:664] <= {8{(wt1_sd_nz[83] | wt1_sd_nan[41])}} & wt1_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[679:672] <= {8{(wt1_sd_nz[84] | wt1_sd_nan[42])}} & wt1_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[687:680] <= {8{(wt1_sd_nz[85] | wt1_sd_nan[42])}} & wt1_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[695:688] <= {8{(wt1_sd_nz[86] | wt1_sd_nan[43])}} & wt1_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[703:696] <= {8{(wt1_sd_nz[87] | wt1_sd_nan[43])}} & wt1_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[711:704] <= {8{(wt1_sd_nz[88] | wt1_sd_nan[44])}} & wt1_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[719:712] <= {8{(wt1_sd_nz[89] | wt1_sd_nan[44])}} & wt1_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[727:720] <= {8{(wt1_sd_nz[90] | wt1_sd_nan[45])}} & wt1_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[735:728] <= {8{(wt1_sd_nz[91] | wt1_sd_nan[45])}} & wt1_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[743:736] <= {8{(wt1_sd_nz[92] | wt1_sd_nan[46])}} & wt1_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[751:744] <= {8{(wt1_sd_nz[93] | wt1_sd_nan[46])}} & wt1_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[759:752] <= {8{(wt1_sd_nz[94] | wt1_sd_nan[47])}} & wt1_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[767:760] <= {8{(wt1_sd_nz[95] | wt1_sd_nan[47])}} & wt1_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[775:768] <= {8{(wt1_sd_nz[96] | wt1_sd_nan[48])}} & wt1_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[783:776] <= {8{(wt1_sd_nz[97] | wt1_sd_nan[48])}} & wt1_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[791:784] <= {8{(wt1_sd_nz[98] | wt1_sd_nan[49])}} & wt1_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[799:792] <= {8{(wt1_sd_nz[99] | wt1_sd_nan[49])}} & wt1_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[807:800] <= {8{(wt1_sd_nz[100] | wt1_sd_nan[50])}} & wt1_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[815:808] <= {8{(wt1_sd_nz[101] | wt1_sd_nan[50])}} & wt1_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[823:816] <= {8{(wt1_sd_nz[102] | wt1_sd_nan[51])}} & wt1_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[831:824] <= {8{(wt1_sd_nz[103] | wt1_sd_nan[51])}} & wt1_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[839:832] <= {8{(wt1_sd_nz[104] | wt1_sd_nan[52])}} & wt1_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[847:840] <= {8{(wt1_sd_nz[105] | wt1_sd_nan[52])}} & wt1_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[855:848] <= {8{(wt1_sd_nz[106] | wt1_sd_nan[53])}} & wt1_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[863:856] <= {8{(wt1_sd_nz[107] | wt1_sd_nan[53])}} & wt1_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[871:864] <= {8{(wt1_sd_nz[108] | wt1_sd_nan[54])}} & wt1_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[879:872] <= {8{(wt1_sd_nz[109] | wt1_sd_nan[54])}} & wt1_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[887:880] <= {8{(wt1_sd_nz[110] | wt1_sd_nan[55])}} & wt1_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[895:888] <= {8{(wt1_sd_nz[111] | wt1_sd_nan[55])}} & wt1_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[903:896] <= {8{(wt1_sd_nz[112] | wt1_sd_nan[56])}} & wt1_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[911:904] <= {8{(wt1_sd_nz[113] | wt1_sd_nan[56])}} & wt1_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[919:912] <= {8{(wt1_sd_nz[114] | wt1_sd_nan[57])}} & wt1_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[927:920] <= {8{(wt1_sd_nz[115] | wt1_sd_nan[57])}} & wt1_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[935:928] <= {8{(wt1_sd_nz[116] | wt1_sd_nan[58])}} & wt1_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[943:936] <= {8{(wt1_sd_nz[117] | wt1_sd_nan[58])}} & wt1_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[951:944] <= {8{(wt1_sd_nz[118] | wt1_sd_nan[59])}} & wt1_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[959:952] <= {8{(wt1_sd_nz[119] | wt1_sd_nan[59])}} & wt1_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[967:960] <= {8{(wt1_sd_nz[120] | wt1_sd_nan[60])}} & wt1_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[975:968] <= {8{(wt1_sd_nz[121] | wt1_sd_nan[60])}} & wt1_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[983:976] <= {8{(wt1_sd_nz[122] | wt1_sd_nan[61])}} & wt1_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[991:984] <= {8{(wt1_sd_nz[123] | wt1_sd_nan[61])}} & wt1_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[999:992] <= {8{(wt1_sd_nz[124] | wt1_sd_nan[62])}} & wt1_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[1007:1000] <= {8{(wt1_sd_nz[125] | wt1_sd_nan[62])}} & wt1_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[1015:1008] <= {8{(wt1_sd_nz[126] | wt1_sd_nan[63])}} & wt1_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b1) begin
    wt1_actv_data[1023:1016] <= {8{(wt1_sd_nz[127] | wt1_sd_nan[63])}} & wt1_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[1] & wt1_actv_pvld_w) == 1'b0) begin
  end else begin
    wt1_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt2_sd_pvld
  or dat_actv_stripe_end
  or wt2_actv_vld
  ) begin
    wt2_actv_pvld_w = dat_pre_stripe_st[2] ? wt2_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt2_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt2_actv_vld <= 1'b0;
  end else begin
  wt2_actv_vld <= wt2_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt2_actv_pvld <= {104{1'b0}};
  end else begin
  wt2_actv_pvld <= {104{wt2_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_nz <= wt2_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w & cfg_is_fp16_d1[76]) == 1'b1) begin
    wt2_actv_nan <= wt2_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w & cfg_is_fp16_d1[76]) == 1'b0) begin
  end else begin
    wt2_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[7:0] <= {8{(wt2_sd_nz[0] | wt2_sd_nan[0])}} & wt2_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[15:8] <= {8{(wt2_sd_nz[1] | wt2_sd_nan[0])}} & wt2_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[23:16] <= {8{(wt2_sd_nz[2] | wt2_sd_nan[1])}} & wt2_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[31:24] <= {8{(wt2_sd_nz[3] | wt2_sd_nan[1])}} & wt2_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[39:32] <= {8{(wt2_sd_nz[4] | wt2_sd_nan[2])}} & wt2_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[47:40] <= {8{(wt2_sd_nz[5] | wt2_sd_nan[2])}} & wt2_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[55:48] <= {8{(wt2_sd_nz[6] | wt2_sd_nan[3])}} & wt2_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[63:56] <= {8{(wt2_sd_nz[7] | wt2_sd_nan[3])}} & wt2_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[71:64] <= {8{(wt2_sd_nz[8] | wt2_sd_nan[4])}} & wt2_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[79:72] <= {8{(wt2_sd_nz[9] | wt2_sd_nan[4])}} & wt2_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[87:80] <= {8{(wt2_sd_nz[10] | wt2_sd_nan[5])}} & wt2_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[95:88] <= {8{(wt2_sd_nz[11] | wt2_sd_nan[5])}} & wt2_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[103:96] <= {8{(wt2_sd_nz[12] | wt2_sd_nan[6])}} & wt2_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[111:104] <= {8{(wt2_sd_nz[13] | wt2_sd_nan[6])}} & wt2_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[119:112] <= {8{(wt2_sd_nz[14] | wt2_sd_nan[7])}} & wt2_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[127:120] <= {8{(wt2_sd_nz[15] | wt2_sd_nan[7])}} & wt2_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[135:128] <= {8{(wt2_sd_nz[16] | wt2_sd_nan[8])}} & wt2_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[143:136] <= {8{(wt2_sd_nz[17] | wt2_sd_nan[8])}} & wt2_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[151:144] <= {8{(wt2_sd_nz[18] | wt2_sd_nan[9])}} & wt2_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[159:152] <= {8{(wt2_sd_nz[19] | wt2_sd_nan[9])}} & wt2_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[167:160] <= {8{(wt2_sd_nz[20] | wt2_sd_nan[10])}} & wt2_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[175:168] <= {8{(wt2_sd_nz[21] | wt2_sd_nan[10])}} & wt2_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[183:176] <= {8{(wt2_sd_nz[22] | wt2_sd_nan[11])}} & wt2_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[191:184] <= {8{(wt2_sd_nz[23] | wt2_sd_nan[11])}} & wt2_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[199:192] <= {8{(wt2_sd_nz[24] | wt2_sd_nan[12])}} & wt2_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[207:200] <= {8{(wt2_sd_nz[25] | wt2_sd_nan[12])}} & wt2_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[215:208] <= {8{(wt2_sd_nz[26] | wt2_sd_nan[13])}} & wt2_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[223:216] <= {8{(wt2_sd_nz[27] | wt2_sd_nan[13])}} & wt2_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[231:224] <= {8{(wt2_sd_nz[28] | wt2_sd_nan[14])}} & wt2_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[239:232] <= {8{(wt2_sd_nz[29] | wt2_sd_nan[14])}} & wt2_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[247:240] <= {8{(wt2_sd_nz[30] | wt2_sd_nan[15])}} & wt2_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[255:248] <= {8{(wt2_sd_nz[31] | wt2_sd_nan[15])}} & wt2_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[263:256] <= {8{(wt2_sd_nz[32] | wt2_sd_nan[16])}} & wt2_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[271:264] <= {8{(wt2_sd_nz[33] | wt2_sd_nan[16])}} & wt2_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[279:272] <= {8{(wt2_sd_nz[34] | wt2_sd_nan[17])}} & wt2_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[287:280] <= {8{(wt2_sd_nz[35] | wt2_sd_nan[17])}} & wt2_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[295:288] <= {8{(wt2_sd_nz[36] | wt2_sd_nan[18])}} & wt2_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[303:296] <= {8{(wt2_sd_nz[37] | wt2_sd_nan[18])}} & wt2_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[311:304] <= {8{(wt2_sd_nz[38] | wt2_sd_nan[19])}} & wt2_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[319:312] <= {8{(wt2_sd_nz[39] | wt2_sd_nan[19])}} & wt2_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[327:320] <= {8{(wt2_sd_nz[40] | wt2_sd_nan[20])}} & wt2_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[335:328] <= {8{(wt2_sd_nz[41] | wt2_sd_nan[20])}} & wt2_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[343:336] <= {8{(wt2_sd_nz[42] | wt2_sd_nan[21])}} & wt2_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[351:344] <= {8{(wt2_sd_nz[43] | wt2_sd_nan[21])}} & wt2_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[359:352] <= {8{(wt2_sd_nz[44] | wt2_sd_nan[22])}} & wt2_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[367:360] <= {8{(wt2_sd_nz[45] | wt2_sd_nan[22])}} & wt2_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[375:368] <= {8{(wt2_sd_nz[46] | wt2_sd_nan[23])}} & wt2_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[383:376] <= {8{(wt2_sd_nz[47] | wt2_sd_nan[23])}} & wt2_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[391:384] <= {8{(wt2_sd_nz[48] | wt2_sd_nan[24])}} & wt2_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[399:392] <= {8{(wt2_sd_nz[49] | wt2_sd_nan[24])}} & wt2_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[407:400] <= {8{(wt2_sd_nz[50] | wt2_sd_nan[25])}} & wt2_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[415:408] <= {8{(wt2_sd_nz[51] | wt2_sd_nan[25])}} & wt2_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[423:416] <= {8{(wt2_sd_nz[52] | wt2_sd_nan[26])}} & wt2_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[431:424] <= {8{(wt2_sd_nz[53] | wt2_sd_nan[26])}} & wt2_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[439:432] <= {8{(wt2_sd_nz[54] | wt2_sd_nan[27])}} & wt2_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[447:440] <= {8{(wt2_sd_nz[55] | wt2_sd_nan[27])}} & wt2_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[455:448] <= {8{(wt2_sd_nz[56] | wt2_sd_nan[28])}} & wt2_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[463:456] <= {8{(wt2_sd_nz[57] | wt2_sd_nan[28])}} & wt2_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[471:464] <= {8{(wt2_sd_nz[58] | wt2_sd_nan[29])}} & wt2_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[479:472] <= {8{(wt2_sd_nz[59] | wt2_sd_nan[29])}} & wt2_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[487:480] <= {8{(wt2_sd_nz[60] | wt2_sd_nan[30])}} & wt2_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[495:488] <= {8{(wt2_sd_nz[61] | wt2_sd_nan[30])}} & wt2_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[503:496] <= {8{(wt2_sd_nz[62] | wt2_sd_nan[31])}} & wt2_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[511:504] <= {8{(wt2_sd_nz[63] | wt2_sd_nan[31])}} & wt2_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[519:512] <= {8{(wt2_sd_nz[64] | wt2_sd_nan[32])}} & wt2_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[527:520] <= {8{(wt2_sd_nz[65] | wt2_sd_nan[32])}} & wt2_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[535:528] <= {8{(wt2_sd_nz[66] | wt2_sd_nan[33])}} & wt2_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[543:536] <= {8{(wt2_sd_nz[67] | wt2_sd_nan[33])}} & wt2_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[551:544] <= {8{(wt2_sd_nz[68] | wt2_sd_nan[34])}} & wt2_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[559:552] <= {8{(wt2_sd_nz[69] | wt2_sd_nan[34])}} & wt2_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[567:560] <= {8{(wt2_sd_nz[70] | wt2_sd_nan[35])}} & wt2_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[575:568] <= {8{(wt2_sd_nz[71] | wt2_sd_nan[35])}} & wt2_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[583:576] <= {8{(wt2_sd_nz[72] | wt2_sd_nan[36])}} & wt2_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[591:584] <= {8{(wt2_sd_nz[73] | wt2_sd_nan[36])}} & wt2_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[599:592] <= {8{(wt2_sd_nz[74] | wt2_sd_nan[37])}} & wt2_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[607:600] <= {8{(wt2_sd_nz[75] | wt2_sd_nan[37])}} & wt2_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[615:608] <= {8{(wt2_sd_nz[76] | wt2_sd_nan[38])}} & wt2_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[623:616] <= {8{(wt2_sd_nz[77] | wt2_sd_nan[38])}} & wt2_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[631:624] <= {8{(wt2_sd_nz[78] | wt2_sd_nan[39])}} & wt2_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[639:632] <= {8{(wt2_sd_nz[79] | wt2_sd_nan[39])}} & wt2_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[647:640] <= {8{(wt2_sd_nz[80] | wt2_sd_nan[40])}} & wt2_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[655:648] <= {8{(wt2_sd_nz[81] | wt2_sd_nan[40])}} & wt2_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[663:656] <= {8{(wt2_sd_nz[82] | wt2_sd_nan[41])}} & wt2_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[671:664] <= {8{(wt2_sd_nz[83] | wt2_sd_nan[41])}} & wt2_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[679:672] <= {8{(wt2_sd_nz[84] | wt2_sd_nan[42])}} & wt2_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[687:680] <= {8{(wt2_sd_nz[85] | wt2_sd_nan[42])}} & wt2_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[695:688] <= {8{(wt2_sd_nz[86] | wt2_sd_nan[43])}} & wt2_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[703:696] <= {8{(wt2_sd_nz[87] | wt2_sd_nan[43])}} & wt2_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[711:704] <= {8{(wt2_sd_nz[88] | wt2_sd_nan[44])}} & wt2_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[719:712] <= {8{(wt2_sd_nz[89] | wt2_sd_nan[44])}} & wt2_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[727:720] <= {8{(wt2_sd_nz[90] | wt2_sd_nan[45])}} & wt2_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[735:728] <= {8{(wt2_sd_nz[91] | wt2_sd_nan[45])}} & wt2_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[743:736] <= {8{(wt2_sd_nz[92] | wt2_sd_nan[46])}} & wt2_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[751:744] <= {8{(wt2_sd_nz[93] | wt2_sd_nan[46])}} & wt2_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[759:752] <= {8{(wt2_sd_nz[94] | wt2_sd_nan[47])}} & wt2_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[767:760] <= {8{(wt2_sd_nz[95] | wt2_sd_nan[47])}} & wt2_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[775:768] <= {8{(wt2_sd_nz[96] | wt2_sd_nan[48])}} & wt2_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[783:776] <= {8{(wt2_sd_nz[97] | wt2_sd_nan[48])}} & wt2_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[791:784] <= {8{(wt2_sd_nz[98] | wt2_sd_nan[49])}} & wt2_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[799:792] <= {8{(wt2_sd_nz[99] | wt2_sd_nan[49])}} & wt2_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[807:800] <= {8{(wt2_sd_nz[100] | wt2_sd_nan[50])}} & wt2_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[815:808] <= {8{(wt2_sd_nz[101] | wt2_sd_nan[50])}} & wt2_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[823:816] <= {8{(wt2_sd_nz[102] | wt2_sd_nan[51])}} & wt2_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[831:824] <= {8{(wt2_sd_nz[103] | wt2_sd_nan[51])}} & wt2_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[839:832] <= {8{(wt2_sd_nz[104] | wt2_sd_nan[52])}} & wt2_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[847:840] <= {8{(wt2_sd_nz[105] | wt2_sd_nan[52])}} & wt2_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[855:848] <= {8{(wt2_sd_nz[106] | wt2_sd_nan[53])}} & wt2_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[863:856] <= {8{(wt2_sd_nz[107] | wt2_sd_nan[53])}} & wt2_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[871:864] <= {8{(wt2_sd_nz[108] | wt2_sd_nan[54])}} & wt2_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[879:872] <= {8{(wt2_sd_nz[109] | wt2_sd_nan[54])}} & wt2_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[887:880] <= {8{(wt2_sd_nz[110] | wt2_sd_nan[55])}} & wt2_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[895:888] <= {8{(wt2_sd_nz[111] | wt2_sd_nan[55])}} & wt2_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[903:896] <= {8{(wt2_sd_nz[112] | wt2_sd_nan[56])}} & wt2_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[911:904] <= {8{(wt2_sd_nz[113] | wt2_sd_nan[56])}} & wt2_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[919:912] <= {8{(wt2_sd_nz[114] | wt2_sd_nan[57])}} & wt2_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[927:920] <= {8{(wt2_sd_nz[115] | wt2_sd_nan[57])}} & wt2_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[935:928] <= {8{(wt2_sd_nz[116] | wt2_sd_nan[58])}} & wt2_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[943:936] <= {8{(wt2_sd_nz[117] | wt2_sd_nan[58])}} & wt2_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[951:944] <= {8{(wt2_sd_nz[118] | wt2_sd_nan[59])}} & wt2_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[959:952] <= {8{(wt2_sd_nz[119] | wt2_sd_nan[59])}} & wt2_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[967:960] <= {8{(wt2_sd_nz[120] | wt2_sd_nan[60])}} & wt2_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[975:968] <= {8{(wt2_sd_nz[121] | wt2_sd_nan[60])}} & wt2_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[983:976] <= {8{(wt2_sd_nz[122] | wt2_sd_nan[61])}} & wt2_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[991:984] <= {8{(wt2_sd_nz[123] | wt2_sd_nan[61])}} & wt2_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[999:992] <= {8{(wt2_sd_nz[124] | wt2_sd_nan[62])}} & wt2_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[1007:1000] <= {8{(wt2_sd_nz[125] | wt2_sd_nan[62])}} & wt2_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[1015:1008] <= {8{(wt2_sd_nz[126] | wt2_sd_nan[63])}} & wt2_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b1) begin
    wt2_actv_data[1023:1016] <= {8{(wt2_sd_nz[127] | wt2_sd_nan[63])}} & wt2_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[2] & wt2_actv_pvld_w) == 1'b0) begin
  end else begin
    wt2_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt3_sd_pvld
  or dat_actv_stripe_end
  or wt3_actv_vld
  ) begin
    wt3_actv_pvld_w = dat_pre_stripe_st[3] ? wt3_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt3_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt3_actv_vld <= 1'b0;
  end else begin
  wt3_actv_vld <= wt3_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt3_actv_pvld <= {104{1'b0}};
  end else begin
  wt3_actv_pvld <= {104{wt3_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_nz <= wt3_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w & cfg_is_fp16_d1[77]) == 1'b1) begin
    wt3_actv_nan <= wt3_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w & cfg_is_fp16_d1[77]) == 1'b0) begin
  end else begin
    wt3_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[7:0] <= {8{(wt3_sd_nz[0] | wt3_sd_nan[0])}} & wt3_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[15:8] <= {8{(wt3_sd_nz[1] | wt3_sd_nan[0])}} & wt3_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[23:16] <= {8{(wt3_sd_nz[2] | wt3_sd_nan[1])}} & wt3_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[31:24] <= {8{(wt3_sd_nz[3] | wt3_sd_nan[1])}} & wt3_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[39:32] <= {8{(wt3_sd_nz[4] | wt3_sd_nan[2])}} & wt3_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[47:40] <= {8{(wt3_sd_nz[5] | wt3_sd_nan[2])}} & wt3_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[55:48] <= {8{(wt3_sd_nz[6] | wt3_sd_nan[3])}} & wt3_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[63:56] <= {8{(wt3_sd_nz[7] | wt3_sd_nan[3])}} & wt3_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[71:64] <= {8{(wt3_sd_nz[8] | wt3_sd_nan[4])}} & wt3_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[79:72] <= {8{(wt3_sd_nz[9] | wt3_sd_nan[4])}} & wt3_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[87:80] <= {8{(wt3_sd_nz[10] | wt3_sd_nan[5])}} & wt3_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[95:88] <= {8{(wt3_sd_nz[11] | wt3_sd_nan[5])}} & wt3_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[103:96] <= {8{(wt3_sd_nz[12] | wt3_sd_nan[6])}} & wt3_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[111:104] <= {8{(wt3_sd_nz[13] | wt3_sd_nan[6])}} & wt3_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[119:112] <= {8{(wt3_sd_nz[14] | wt3_sd_nan[7])}} & wt3_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[127:120] <= {8{(wt3_sd_nz[15] | wt3_sd_nan[7])}} & wt3_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[135:128] <= {8{(wt3_sd_nz[16] | wt3_sd_nan[8])}} & wt3_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[143:136] <= {8{(wt3_sd_nz[17] | wt3_sd_nan[8])}} & wt3_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[151:144] <= {8{(wt3_sd_nz[18] | wt3_sd_nan[9])}} & wt3_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[159:152] <= {8{(wt3_sd_nz[19] | wt3_sd_nan[9])}} & wt3_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[167:160] <= {8{(wt3_sd_nz[20] | wt3_sd_nan[10])}} & wt3_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[175:168] <= {8{(wt3_sd_nz[21] | wt3_sd_nan[10])}} & wt3_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[183:176] <= {8{(wt3_sd_nz[22] | wt3_sd_nan[11])}} & wt3_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[191:184] <= {8{(wt3_sd_nz[23] | wt3_sd_nan[11])}} & wt3_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[199:192] <= {8{(wt3_sd_nz[24] | wt3_sd_nan[12])}} & wt3_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[207:200] <= {8{(wt3_sd_nz[25] | wt3_sd_nan[12])}} & wt3_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[215:208] <= {8{(wt3_sd_nz[26] | wt3_sd_nan[13])}} & wt3_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[223:216] <= {8{(wt3_sd_nz[27] | wt3_sd_nan[13])}} & wt3_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[231:224] <= {8{(wt3_sd_nz[28] | wt3_sd_nan[14])}} & wt3_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[239:232] <= {8{(wt3_sd_nz[29] | wt3_sd_nan[14])}} & wt3_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[247:240] <= {8{(wt3_sd_nz[30] | wt3_sd_nan[15])}} & wt3_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[255:248] <= {8{(wt3_sd_nz[31] | wt3_sd_nan[15])}} & wt3_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[263:256] <= {8{(wt3_sd_nz[32] | wt3_sd_nan[16])}} & wt3_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[271:264] <= {8{(wt3_sd_nz[33] | wt3_sd_nan[16])}} & wt3_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[279:272] <= {8{(wt3_sd_nz[34] | wt3_sd_nan[17])}} & wt3_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[287:280] <= {8{(wt3_sd_nz[35] | wt3_sd_nan[17])}} & wt3_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[295:288] <= {8{(wt3_sd_nz[36] | wt3_sd_nan[18])}} & wt3_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[303:296] <= {8{(wt3_sd_nz[37] | wt3_sd_nan[18])}} & wt3_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[311:304] <= {8{(wt3_sd_nz[38] | wt3_sd_nan[19])}} & wt3_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[319:312] <= {8{(wt3_sd_nz[39] | wt3_sd_nan[19])}} & wt3_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[327:320] <= {8{(wt3_sd_nz[40] | wt3_sd_nan[20])}} & wt3_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[335:328] <= {8{(wt3_sd_nz[41] | wt3_sd_nan[20])}} & wt3_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[343:336] <= {8{(wt3_sd_nz[42] | wt3_sd_nan[21])}} & wt3_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[351:344] <= {8{(wt3_sd_nz[43] | wt3_sd_nan[21])}} & wt3_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[359:352] <= {8{(wt3_sd_nz[44] | wt3_sd_nan[22])}} & wt3_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[367:360] <= {8{(wt3_sd_nz[45] | wt3_sd_nan[22])}} & wt3_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[375:368] <= {8{(wt3_sd_nz[46] | wt3_sd_nan[23])}} & wt3_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[383:376] <= {8{(wt3_sd_nz[47] | wt3_sd_nan[23])}} & wt3_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[391:384] <= {8{(wt3_sd_nz[48] | wt3_sd_nan[24])}} & wt3_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[399:392] <= {8{(wt3_sd_nz[49] | wt3_sd_nan[24])}} & wt3_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[407:400] <= {8{(wt3_sd_nz[50] | wt3_sd_nan[25])}} & wt3_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[415:408] <= {8{(wt3_sd_nz[51] | wt3_sd_nan[25])}} & wt3_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[423:416] <= {8{(wt3_sd_nz[52] | wt3_sd_nan[26])}} & wt3_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[431:424] <= {8{(wt3_sd_nz[53] | wt3_sd_nan[26])}} & wt3_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[439:432] <= {8{(wt3_sd_nz[54] | wt3_sd_nan[27])}} & wt3_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[447:440] <= {8{(wt3_sd_nz[55] | wt3_sd_nan[27])}} & wt3_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[455:448] <= {8{(wt3_sd_nz[56] | wt3_sd_nan[28])}} & wt3_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[463:456] <= {8{(wt3_sd_nz[57] | wt3_sd_nan[28])}} & wt3_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[471:464] <= {8{(wt3_sd_nz[58] | wt3_sd_nan[29])}} & wt3_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[479:472] <= {8{(wt3_sd_nz[59] | wt3_sd_nan[29])}} & wt3_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[487:480] <= {8{(wt3_sd_nz[60] | wt3_sd_nan[30])}} & wt3_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[495:488] <= {8{(wt3_sd_nz[61] | wt3_sd_nan[30])}} & wt3_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[503:496] <= {8{(wt3_sd_nz[62] | wt3_sd_nan[31])}} & wt3_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[511:504] <= {8{(wt3_sd_nz[63] | wt3_sd_nan[31])}} & wt3_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[519:512] <= {8{(wt3_sd_nz[64] | wt3_sd_nan[32])}} & wt3_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[527:520] <= {8{(wt3_sd_nz[65] | wt3_sd_nan[32])}} & wt3_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[535:528] <= {8{(wt3_sd_nz[66] | wt3_sd_nan[33])}} & wt3_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[543:536] <= {8{(wt3_sd_nz[67] | wt3_sd_nan[33])}} & wt3_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[551:544] <= {8{(wt3_sd_nz[68] | wt3_sd_nan[34])}} & wt3_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[559:552] <= {8{(wt3_sd_nz[69] | wt3_sd_nan[34])}} & wt3_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[567:560] <= {8{(wt3_sd_nz[70] | wt3_sd_nan[35])}} & wt3_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[575:568] <= {8{(wt3_sd_nz[71] | wt3_sd_nan[35])}} & wt3_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[583:576] <= {8{(wt3_sd_nz[72] | wt3_sd_nan[36])}} & wt3_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[591:584] <= {8{(wt3_sd_nz[73] | wt3_sd_nan[36])}} & wt3_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[599:592] <= {8{(wt3_sd_nz[74] | wt3_sd_nan[37])}} & wt3_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[607:600] <= {8{(wt3_sd_nz[75] | wt3_sd_nan[37])}} & wt3_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[615:608] <= {8{(wt3_sd_nz[76] | wt3_sd_nan[38])}} & wt3_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[623:616] <= {8{(wt3_sd_nz[77] | wt3_sd_nan[38])}} & wt3_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[631:624] <= {8{(wt3_sd_nz[78] | wt3_sd_nan[39])}} & wt3_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[639:632] <= {8{(wt3_sd_nz[79] | wt3_sd_nan[39])}} & wt3_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[647:640] <= {8{(wt3_sd_nz[80] | wt3_sd_nan[40])}} & wt3_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[655:648] <= {8{(wt3_sd_nz[81] | wt3_sd_nan[40])}} & wt3_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[663:656] <= {8{(wt3_sd_nz[82] | wt3_sd_nan[41])}} & wt3_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[671:664] <= {8{(wt3_sd_nz[83] | wt3_sd_nan[41])}} & wt3_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[679:672] <= {8{(wt3_sd_nz[84] | wt3_sd_nan[42])}} & wt3_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[687:680] <= {8{(wt3_sd_nz[85] | wt3_sd_nan[42])}} & wt3_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[695:688] <= {8{(wt3_sd_nz[86] | wt3_sd_nan[43])}} & wt3_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[703:696] <= {8{(wt3_sd_nz[87] | wt3_sd_nan[43])}} & wt3_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[711:704] <= {8{(wt3_sd_nz[88] | wt3_sd_nan[44])}} & wt3_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[719:712] <= {8{(wt3_sd_nz[89] | wt3_sd_nan[44])}} & wt3_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[727:720] <= {8{(wt3_sd_nz[90] | wt3_sd_nan[45])}} & wt3_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[735:728] <= {8{(wt3_sd_nz[91] | wt3_sd_nan[45])}} & wt3_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[743:736] <= {8{(wt3_sd_nz[92] | wt3_sd_nan[46])}} & wt3_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[751:744] <= {8{(wt3_sd_nz[93] | wt3_sd_nan[46])}} & wt3_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[759:752] <= {8{(wt3_sd_nz[94] | wt3_sd_nan[47])}} & wt3_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[767:760] <= {8{(wt3_sd_nz[95] | wt3_sd_nan[47])}} & wt3_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[775:768] <= {8{(wt3_sd_nz[96] | wt3_sd_nan[48])}} & wt3_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[783:776] <= {8{(wt3_sd_nz[97] | wt3_sd_nan[48])}} & wt3_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[791:784] <= {8{(wt3_sd_nz[98] | wt3_sd_nan[49])}} & wt3_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[799:792] <= {8{(wt3_sd_nz[99] | wt3_sd_nan[49])}} & wt3_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[807:800] <= {8{(wt3_sd_nz[100] | wt3_sd_nan[50])}} & wt3_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[815:808] <= {8{(wt3_sd_nz[101] | wt3_sd_nan[50])}} & wt3_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[823:816] <= {8{(wt3_sd_nz[102] | wt3_sd_nan[51])}} & wt3_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[831:824] <= {8{(wt3_sd_nz[103] | wt3_sd_nan[51])}} & wt3_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[839:832] <= {8{(wt3_sd_nz[104] | wt3_sd_nan[52])}} & wt3_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[847:840] <= {8{(wt3_sd_nz[105] | wt3_sd_nan[52])}} & wt3_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[855:848] <= {8{(wt3_sd_nz[106] | wt3_sd_nan[53])}} & wt3_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[863:856] <= {8{(wt3_sd_nz[107] | wt3_sd_nan[53])}} & wt3_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[871:864] <= {8{(wt3_sd_nz[108] | wt3_sd_nan[54])}} & wt3_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[879:872] <= {8{(wt3_sd_nz[109] | wt3_sd_nan[54])}} & wt3_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[887:880] <= {8{(wt3_sd_nz[110] | wt3_sd_nan[55])}} & wt3_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[895:888] <= {8{(wt3_sd_nz[111] | wt3_sd_nan[55])}} & wt3_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[903:896] <= {8{(wt3_sd_nz[112] | wt3_sd_nan[56])}} & wt3_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[911:904] <= {8{(wt3_sd_nz[113] | wt3_sd_nan[56])}} & wt3_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[919:912] <= {8{(wt3_sd_nz[114] | wt3_sd_nan[57])}} & wt3_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[927:920] <= {8{(wt3_sd_nz[115] | wt3_sd_nan[57])}} & wt3_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[935:928] <= {8{(wt3_sd_nz[116] | wt3_sd_nan[58])}} & wt3_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[943:936] <= {8{(wt3_sd_nz[117] | wt3_sd_nan[58])}} & wt3_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[951:944] <= {8{(wt3_sd_nz[118] | wt3_sd_nan[59])}} & wt3_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[959:952] <= {8{(wt3_sd_nz[119] | wt3_sd_nan[59])}} & wt3_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[967:960] <= {8{(wt3_sd_nz[120] | wt3_sd_nan[60])}} & wt3_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[975:968] <= {8{(wt3_sd_nz[121] | wt3_sd_nan[60])}} & wt3_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[983:976] <= {8{(wt3_sd_nz[122] | wt3_sd_nan[61])}} & wt3_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[991:984] <= {8{(wt3_sd_nz[123] | wt3_sd_nan[61])}} & wt3_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[999:992] <= {8{(wt3_sd_nz[124] | wt3_sd_nan[62])}} & wt3_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[1007:1000] <= {8{(wt3_sd_nz[125] | wt3_sd_nan[62])}} & wt3_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[1015:1008] <= {8{(wt3_sd_nz[126] | wt3_sd_nan[63])}} & wt3_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b1) begin
    wt3_actv_data[1023:1016] <= {8{(wt3_sd_nz[127] | wt3_sd_nan[63])}} & wt3_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[3] & wt3_actv_pvld_w) == 1'b0) begin
  end else begin
    wt3_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt4_sd_pvld
  or dat_actv_stripe_end
  or wt4_actv_vld
  ) begin
    wt4_actv_pvld_w = dat_pre_stripe_st[4] ? wt4_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt4_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt4_actv_vld <= 1'b0;
  end else begin
  wt4_actv_vld <= wt4_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt4_actv_pvld <= {104{1'b0}};
  end else begin
  wt4_actv_pvld <= {104{wt4_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_nz <= wt4_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w & cfg_is_fp16_d1[78]) == 1'b1) begin
    wt4_actv_nan <= wt4_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w & cfg_is_fp16_d1[78]) == 1'b0) begin
  end else begin
    wt4_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[7:0] <= {8{(wt4_sd_nz[0] | wt4_sd_nan[0])}} & wt4_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[15:8] <= {8{(wt4_sd_nz[1] | wt4_sd_nan[0])}} & wt4_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[23:16] <= {8{(wt4_sd_nz[2] | wt4_sd_nan[1])}} & wt4_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[31:24] <= {8{(wt4_sd_nz[3] | wt4_sd_nan[1])}} & wt4_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[39:32] <= {8{(wt4_sd_nz[4] | wt4_sd_nan[2])}} & wt4_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[47:40] <= {8{(wt4_sd_nz[5] | wt4_sd_nan[2])}} & wt4_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[55:48] <= {8{(wt4_sd_nz[6] | wt4_sd_nan[3])}} & wt4_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[63:56] <= {8{(wt4_sd_nz[7] | wt4_sd_nan[3])}} & wt4_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[71:64] <= {8{(wt4_sd_nz[8] | wt4_sd_nan[4])}} & wt4_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[79:72] <= {8{(wt4_sd_nz[9] | wt4_sd_nan[4])}} & wt4_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[87:80] <= {8{(wt4_sd_nz[10] | wt4_sd_nan[5])}} & wt4_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[95:88] <= {8{(wt4_sd_nz[11] | wt4_sd_nan[5])}} & wt4_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[103:96] <= {8{(wt4_sd_nz[12] | wt4_sd_nan[6])}} & wt4_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[111:104] <= {8{(wt4_sd_nz[13] | wt4_sd_nan[6])}} & wt4_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[119:112] <= {8{(wt4_sd_nz[14] | wt4_sd_nan[7])}} & wt4_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[127:120] <= {8{(wt4_sd_nz[15] | wt4_sd_nan[7])}} & wt4_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[135:128] <= {8{(wt4_sd_nz[16] | wt4_sd_nan[8])}} & wt4_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[143:136] <= {8{(wt4_sd_nz[17] | wt4_sd_nan[8])}} & wt4_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[151:144] <= {8{(wt4_sd_nz[18] | wt4_sd_nan[9])}} & wt4_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[159:152] <= {8{(wt4_sd_nz[19] | wt4_sd_nan[9])}} & wt4_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[167:160] <= {8{(wt4_sd_nz[20] | wt4_sd_nan[10])}} & wt4_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[175:168] <= {8{(wt4_sd_nz[21] | wt4_sd_nan[10])}} & wt4_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[183:176] <= {8{(wt4_sd_nz[22] | wt4_sd_nan[11])}} & wt4_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[191:184] <= {8{(wt4_sd_nz[23] | wt4_sd_nan[11])}} & wt4_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[199:192] <= {8{(wt4_sd_nz[24] | wt4_sd_nan[12])}} & wt4_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[207:200] <= {8{(wt4_sd_nz[25] | wt4_sd_nan[12])}} & wt4_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[215:208] <= {8{(wt4_sd_nz[26] | wt4_sd_nan[13])}} & wt4_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[223:216] <= {8{(wt4_sd_nz[27] | wt4_sd_nan[13])}} & wt4_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[231:224] <= {8{(wt4_sd_nz[28] | wt4_sd_nan[14])}} & wt4_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[239:232] <= {8{(wt4_sd_nz[29] | wt4_sd_nan[14])}} & wt4_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[247:240] <= {8{(wt4_sd_nz[30] | wt4_sd_nan[15])}} & wt4_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[255:248] <= {8{(wt4_sd_nz[31] | wt4_sd_nan[15])}} & wt4_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[263:256] <= {8{(wt4_sd_nz[32] | wt4_sd_nan[16])}} & wt4_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[271:264] <= {8{(wt4_sd_nz[33] | wt4_sd_nan[16])}} & wt4_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[279:272] <= {8{(wt4_sd_nz[34] | wt4_sd_nan[17])}} & wt4_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[287:280] <= {8{(wt4_sd_nz[35] | wt4_sd_nan[17])}} & wt4_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[295:288] <= {8{(wt4_sd_nz[36] | wt4_sd_nan[18])}} & wt4_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[303:296] <= {8{(wt4_sd_nz[37] | wt4_sd_nan[18])}} & wt4_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[311:304] <= {8{(wt4_sd_nz[38] | wt4_sd_nan[19])}} & wt4_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[319:312] <= {8{(wt4_sd_nz[39] | wt4_sd_nan[19])}} & wt4_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[327:320] <= {8{(wt4_sd_nz[40] | wt4_sd_nan[20])}} & wt4_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[335:328] <= {8{(wt4_sd_nz[41] | wt4_sd_nan[20])}} & wt4_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[343:336] <= {8{(wt4_sd_nz[42] | wt4_sd_nan[21])}} & wt4_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[351:344] <= {8{(wt4_sd_nz[43] | wt4_sd_nan[21])}} & wt4_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[359:352] <= {8{(wt4_sd_nz[44] | wt4_sd_nan[22])}} & wt4_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[367:360] <= {8{(wt4_sd_nz[45] | wt4_sd_nan[22])}} & wt4_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[375:368] <= {8{(wt4_sd_nz[46] | wt4_sd_nan[23])}} & wt4_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[383:376] <= {8{(wt4_sd_nz[47] | wt4_sd_nan[23])}} & wt4_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[391:384] <= {8{(wt4_sd_nz[48] | wt4_sd_nan[24])}} & wt4_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[399:392] <= {8{(wt4_sd_nz[49] | wt4_sd_nan[24])}} & wt4_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[407:400] <= {8{(wt4_sd_nz[50] | wt4_sd_nan[25])}} & wt4_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[415:408] <= {8{(wt4_sd_nz[51] | wt4_sd_nan[25])}} & wt4_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[423:416] <= {8{(wt4_sd_nz[52] | wt4_sd_nan[26])}} & wt4_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[431:424] <= {8{(wt4_sd_nz[53] | wt4_sd_nan[26])}} & wt4_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[439:432] <= {8{(wt4_sd_nz[54] | wt4_sd_nan[27])}} & wt4_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[447:440] <= {8{(wt4_sd_nz[55] | wt4_sd_nan[27])}} & wt4_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[455:448] <= {8{(wt4_sd_nz[56] | wt4_sd_nan[28])}} & wt4_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[463:456] <= {8{(wt4_sd_nz[57] | wt4_sd_nan[28])}} & wt4_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[471:464] <= {8{(wt4_sd_nz[58] | wt4_sd_nan[29])}} & wt4_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[479:472] <= {8{(wt4_sd_nz[59] | wt4_sd_nan[29])}} & wt4_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[487:480] <= {8{(wt4_sd_nz[60] | wt4_sd_nan[30])}} & wt4_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[495:488] <= {8{(wt4_sd_nz[61] | wt4_sd_nan[30])}} & wt4_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[503:496] <= {8{(wt4_sd_nz[62] | wt4_sd_nan[31])}} & wt4_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[511:504] <= {8{(wt4_sd_nz[63] | wt4_sd_nan[31])}} & wt4_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[519:512] <= {8{(wt4_sd_nz[64] | wt4_sd_nan[32])}} & wt4_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[527:520] <= {8{(wt4_sd_nz[65] | wt4_sd_nan[32])}} & wt4_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[535:528] <= {8{(wt4_sd_nz[66] | wt4_sd_nan[33])}} & wt4_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[543:536] <= {8{(wt4_sd_nz[67] | wt4_sd_nan[33])}} & wt4_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[551:544] <= {8{(wt4_sd_nz[68] | wt4_sd_nan[34])}} & wt4_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[559:552] <= {8{(wt4_sd_nz[69] | wt4_sd_nan[34])}} & wt4_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[567:560] <= {8{(wt4_sd_nz[70] | wt4_sd_nan[35])}} & wt4_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[575:568] <= {8{(wt4_sd_nz[71] | wt4_sd_nan[35])}} & wt4_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[583:576] <= {8{(wt4_sd_nz[72] | wt4_sd_nan[36])}} & wt4_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[591:584] <= {8{(wt4_sd_nz[73] | wt4_sd_nan[36])}} & wt4_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[599:592] <= {8{(wt4_sd_nz[74] | wt4_sd_nan[37])}} & wt4_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[607:600] <= {8{(wt4_sd_nz[75] | wt4_sd_nan[37])}} & wt4_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[615:608] <= {8{(wt4_sd_nz[76] | wt4_sd_nan[38])}} & wt4_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[623:616] <= {8{(wt4_sd_nz[77] | wt4_sd_nan[38])}} & wt4_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[631:624] <= {8{(wt4_sd_nz[78] | wt4_sd_nan[39])}} & wt4_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[639:632] <= {8{(wt4_sd_nz[79] | wt4_sd_nan[39])}} & wt4_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[647:640] <= {8{(wt4_sd_nz[80] | wt4_sd_nan[40])}} & wt4_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[655:648] <= {8{(wt4_sd_nz[81] | wt4_sd_nan[40])}} & wt4_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[663:656] <= {8{(wt4_sd_nz[82] | wt4_sd_nan[41])}} & wt4_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[671:664] <= {8{(wt4_sd_nz[83] | wt4_sd_nan[41])}} & wt4_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[679:672] <= {8{(wt4_sd_nz[84] | wt4_sd_nan[42])}} & wt4_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[687:680] <= {8{(wt4_sd_nz[85] | wt4_sd_nan[42])}} & wt4_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[695:688] <= {8{(wt4_sd_nz[86] | wt4_sd_nan[43])}} & wt4_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[703:696] <= {8{(wt4_sd_nz[87] | wt4_sd_nan[43])}} & wt4_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[711:704] <= {8{(wt4_sd_nz[88] | wt4_sd_nan[44])}} & wt4_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[719:712] <= {8{(wt4_sd_nz[89] | wt4_sd_nan[44])}} & wt4_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[727:720] <= {8{(wt4_sd_nz[90] | wt4_sd_nan[45])}} & wt4_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[735:728] <= {8{(wt4_sd_nz[91] | wt4_sd_nan[45])}} & wt4_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[743:736] <= {8{(wt4_sd_nz[92] | wt4_sd_nan[46])}} & wt4_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[751:744] <= {8{(wt4_sd_nz[93] | wt4_sd_nan[46])}} & wt4_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[759:752] <= {8{(wt4_sd_nz[94] | wt4_sd_nan[47])}} & wt4_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[767:760] <= {8{(wt4_sd_nz[95] | wt4_sd_nan[47])}} & wt4_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[775:768] <= {8{(wt4_sd_nz[96] | wt4_sd_nan[48])}} & wt4_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[783:776] <= {8{(wt4_sd_nz[97] | wt4_sd_nan[48])}} & wt4_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[791:784] <= {8{(wt4_sd_nz[98] | wt4_sd_nan[49])}} & wt4_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[799:792] <= {8{(wt4_sd_nz[99] | wt4_sd_nan[49])}} & wt4_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[807:800] <= {8{(wt4_sd_nz[100] | wt4_sd_nan[50])}} & wt4_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[815:808] <= {8{(wt4_sd_nz[101] | wt4_sd_nan[50])}} & wt4_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[823:816] <= {8{(wt4_sd_nz[102] | wt4_sd_nan[51])}} & wt4_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[831:824] <= {8{(wt4_sd_nz[103] | wt4_sd_nan[51])}} & wt4_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[839:832] <= {8{(wt4_sd_nz[104] | wt4_sd_nan[52])}} & wt4_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[847:840] <= {8{(wt4_sd_nz[105] | wt4_sd_nan[52])}} & wt4_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[855:848] <= {8{(wt4_sd_nz[106] | wt4_sd_nan[53])}} & wt4_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[863:856] <= {8{(wt4_sd_nz[107] | wt4_sd_nan[53])}} & wt4_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[871:864] <= {8{(wt4_sd_nz[108] | wt4_sd_nan[54])}} & wt4_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[879:872] <= {8{(wt4_sd_nz[109] | wt4_sd_nan[54])}} & wt4_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[887:880] <= {8{(wt4_sd_nz[110] | wt4_sd_nan[55])}} & wt4_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[895:888] <= {8{(wt4_sd_nz[111] | wt4_sd_nan[55])}} & wt4_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[903:896] <= {8{(wt4_sd_nz[112] | wt4_sd_nan[56])}} & wt4_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[911:904] <= {8{(wt4_sd_nz[113] | wt4_sd_nan[56])}} & wt4_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[919:912] <= {8{(wt4_sd_nz[114] | wt4_sd_nan[57])}} & wt4_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[927:920] <= {8{(wt4_sd_nz[115] | wt4_sd_nan[57])}} & wt4_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[935:928] <= {8{(wt4_sd_nz[116] | wt4_sd_nan[58])}} & wt4_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[943:936] <= {8{(wt4_sd_nz[117] | wt4_sd_nan[58])}} & wt4_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[951:944] <= {8{(wt4_sd_nz[118] | wt4_sd_nan[59])}} & wt4_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[959:952] <= {8{(wt4_sd_nz[119] | wt4_sd_nan[59])}} & wt4_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[967:960] <= {8{(wt4_sd_nz[120] | wt4_sd_nan[60])}} & wt4_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[975:968] <= {8{(wt4_sd_nz[121] | wt4_sd_nan[60])}} & wt4_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[983:976] <= {8{(wt4_sd_nz[122] | wt4_sd_nan[61])}} & wt4_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[991:984] <= {8{(wt4_sd_nz[123] | wt4_sd_nan[61])}} & wt4_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[999:992] <= {8{(wt4_sd_nz[124] | wt4_sd_nan[62])}} & wt4_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[1007:1000] <= {8{(wt4_sd_nz[125] | wt4_sd_nan[62])}} & wt4_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[1015:1008] <= {8{(wt4_sd_nz[126] | wt4_sd_nan[63])}} & wt4_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b1) begin
    wt4_actv_data[1023:1016] <= {8{(wt4_sd_nz[127] | wt4_sd_nan[63])}} & wt4_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[4] & wt4_actv_pvld_w) == 1'b0) begin
  end else begin
    wt4_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt5_sd_pvld
  or dat_actv_stripe_end
  or wt5_actv_vld
  ) begin
    wt5_actv_pvld_w = dat_pre_stripe_st[5] ? wt5_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt5_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt5_actv_vld <= 1'b0;
  end else begin
  wt5_actv_vld <= wt5_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt5_actv_pvld <= {104{1'b0}};
  end else begin
  wt5_actv_pvld <= {104{wt5_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_nz <= wt5_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w & cfg_is_fp16_d1[79]) == 1'b1) begin
    wt5_actv_nan <= wt5_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w & cfg_is_fp16_d1[79]) == 1'b0) begin
  end else begin
    wt5_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[7:0] <= {8{(wt5_sd_nz[0] | wt5_sd_nan[0])}} & wt5_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[15:8] <= {8{(wt5_sd_nz[1] | wt5_sd_nan[0])}} & wt5_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[23:16] <= {8{(wt5_sd_nz[2] | wt5_sd_nan[1])}} & wt5_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[31:24] <= {8{(wt5_sd_nz[3] | wt5_sd_nan[1])}} & wt5_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[39:32] <= {8{(wt5_sd_nz[4] | wt5_sd_nan[2])}} & wt5_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[47:40] <= {8{(wt5_sd_nz[5] | wt5_sd_nan[2])}} & wt5_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[55:48] <= {8{(wt5_sd_nz[6] | wt5_sd_nan[3])}} & wt5_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[63:56] <= {8{(wt5_sd_nz[7] | wt5_sd_nan[3])}} & wt5_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[71:64] <= {8{(wt5_sd_nz[8] | wt5_sd_nan[4])}} & wt5_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[79:72] <= {8{(wt5_sd_nz[9] | wt5_sd_nan[4])}} & wt5_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[87:80] <= {8{(wt5_sd_nz[10] | wt5_sd_nan[5])}} & wt5_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[95:88] <= {8{(wt5_sd_nz[11] | wt5_sd_nan[5])}} & wt5_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[103:96] <= {8{(wt5_sd_nz[12] | wt5_sd_nan[6])}} & wt5_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[111:104] <= {8{(wt5_sd_nz[13] | wt5_sd_nan[6])}} & wt5_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[119:112] <= {8{(wt5_sd_nz[14] | wt5_sd_nan[7])}} & wt5_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[127:120] <= {8{(wt5_sd_nz[15] | wt5_sd_nan[7])}} & wt5_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[135:128] <= {8{(wt5_sd_nz[16] | wt5_sd_nan[8])}} & wt5_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[143:136] <= {8{(wt5_sd_nz[17] | wt5_sd_nan[8])}} & wt5_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[151:144] <= {8{(wt5_sd_nz[18] | wt5_sd_nan[9])}} & wt5_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[159:152] <= {8{(wt5_sd_nz[19] | wt5_sd_nan[9])}} & wt5_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[167:160] <= {8{(wt5_sd_nz[20] | wt5_sd_nan[10])}} & wt5_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[175:168] <= {8{(wt5_sd_nz[21] | wt5_sd_nan[10])}} & wt5_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[183:176] <= {8{(wt5_sd_nz[22] | wt5_sd_nan[11])}} & wt5_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[191:184] <= {8{(wt5_sd_nz[23] | wt5_sd_nan[11])}} & wt5_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[199:192] <= {8{(wt5_sd_nz[24] | wt5_sd_nan[12])}} & wt5_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[207:200] <= {8{(wt5_sd_nz[25] | wt5_sd_nan[12])}} & wt5_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[215:208] <= {8{(wt5_sd_nz[26] | wt5_sd_nan[13])}} & wt5_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[223:216] <= {8{(wt5_sd_nz[27] | wt5_sd_nan[13])}} & wt5_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[231:224] <= {8{(wt5_sd_nz[28] | wt5_sd_nan[14])}} & wt5_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[239:232] <= {8{(wt5_sd_nz[29] | wt5_sd_nan[14])}} & wt5_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[247:240] <= {8{(wt5_sd_nz[30] | wt5_sd_nan[15])}} & wt5_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[255:248] <= {8{(wt5_sd_nz[31] | wt5_sd_nan[15])}} & wt5_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[263:256] <= {8{(wt5_sd_nz[32] | wt5_sd_nan[16])}} & wt5_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[271:264] <= {8{(wt5_sd_nz[33] | wt5_sd_nan[16])}} & wt5_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[279:272] <= {8{(wt5_sd_nz[34] | wt5_sd_nan[17])}} & wt5_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[287:280] <= {8{(wt5_sd_nz[35] | wt5_sd_nan[17])}} & wt5_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[295:288] <= {8{(wt5_sd_nz[36] | wt5_sd_nan[18])}} & wt5_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[303:296] <= {8{(wt5_sd_nz[37] | wt5_sd_nan[18])}} & wt5_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[311:304] <= {8{(wt5_sd_nz[38] | wt5_sd_nan[19])}} & wt5_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[319:312] <= {8{(wt5_sd_nz[39] | wt5_sd_nan[19])}} & wt5_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[327:320] <= {8{(wt5_sd_nz[40] | wt5_sd_nan[20])}} & wt5_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[335:328] <= {8{(wt5_sd_nz[41] | wt5_sd_nan[20])}} & wt5_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[343:336] <= {8{(wt5_sd_nz[42] | wt5_sd_nan[21])}} & wt5_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[351:344] <= {8{(wt5_sd_nz[43] | wt5_sd_nan[21])}} & wt5_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[359:352] <= {8{(wt5_sd_nz[44] | wt5_sd_nan[22])}} & wt5_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[367:360] <= {8{(wt5_sd_nz[45] | wt5_sd_nan[22])}} & wt5_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[375:368] <= {8{(wt5_sd_nz[46] | wt5_sd_nan[23])}} & wt5_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[383:376] <= {8{(wt5_sd_nz[47] | wt5_sd_nan[23])}} & wt5_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[391:384] <= {8{(wt5_sd_nz[48] | wt5_sd_nan[24])}} & wt5_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[399:392] <= {8{(wt5_sd_nz[49] | wt5_sd_nan[24])}} & wt5_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[407:400] <= {8{(wt5_sd_nz[50] | wt5_sd_nan[25])}} & wt5_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[415:408] <= {8{(wt5_sd_nz[51] | wt5_sd_nan[25])}} & wt5_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[423:416] <= {8{(wt5_sd_nz[52] | wt5_sd_nan[26])}} & wt5_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[431:424] <= {8{(wt5_sd_nz[53] | wt5_sd_nan[26])}} & wt5_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[439:432] <= {8{(wt5_sd_nz[54] | wt5_sd_nan[27])}} & wt5_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[447:440] <= {8{(wt5_sd_nz[55] | wt5_sd_nan[27])}} & wt5_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[455:448] <= {8{(wt5_sd_nz[56] | wt5_sd_nan[28])}} & wt5_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[463:456] <= {8{(wt5_sd_nz[57] | wt5_sd_nan[28])}} & wt5_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[471:464] <= {8{(wt5_sd_nz[58] | wt5_sd_nan[29])}} & wt5_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[479:472] <= {8{(wt5_sd_nz[59] | wt5_sd_nan[29])}} & wt5_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[487:480] <= {8{(wt5_sd_nz[60] | wt5_sd_nan[30])}} & wt5_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[495:488] <= {8{(wt5_sd_nz[61] | wt5_sd_nan[30])}} & wt5_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[503:496] <= {8{(wt5_sd_nz[62] | wt5_sd_nan[31])}} & wt5_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[511:504] <= {8{(wt5_sd_nz[63] | wt5_sd_nan[31])}} & wt5_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[519:512] <= {8{(wt5_sd_nz[64] | wt5_sd_nan[32])}} & wt5_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[527:520] <= {8{(wt5_sd_nz[65] | wt5_sd_nan[32])}} & wt5_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[535:528] <= {8{(wt5_sd_nz[66] | wt5_sd_nan[33])}} & wt5_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[543:536] <= {8{(wt5_sd_nz[67] | wt5_sd_nan[33])}} & wt5_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[551:544] <= {8{(wt5_sd_nz[68] | wt5_sd_nan[34])}} & wt5_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[559:552] <= {8{(wt5_sd_nz[69] | wt5_sd_nan[34])}} & wt5_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[567:560] <= {8{(wt5_sd_nz[70] | wt5_sd_nan[35])}} & wt5_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[575:568] <= {8{(wt5_sd_nz[71] | wt5_sd_nan[35])}} & wt5_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[583:576] <= {8{(wt5_sd_nz[72] | wt5_sd_nan[36])}} & wt5_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[591:584] <= {8{(wt5_sd_nz[73] | wt5_sd_nan[36])}} & wt5_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[599:592] <= {8{(wt5_sd_nz[74] | wt5_sd_nan[37])}} & wt5_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[607:600] <= {8{(wt5_sd_nz[75] | wt5_sd_nan[37])}} & wt5_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[615:608] <= {8{(wt5_sd_nz[76] | wt5_sd_nan[38])}} & wt5_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[623:616] <= {8{(wt5_sd_nz[77] | wt5_sd_nan[38])}} & wt5_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[631:624] <= {8{(wt5_sd_nz[78] | wt5_sd_nan[39])}} & wt5_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[639:632] <= {8{(wt5_sd_nz[79] | wt5_sd_nan[39])}} & wt5_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[647:640] <= {8{(wt5_sd_nz[80] | wt5_sd_nan[40])}} & wt5_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[655:648] <= {8{(wt5_sd_nz[81] | wt5_sd_nan[40])}} & wt5_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[663:656] <= {8{(wt5_sd_nz[82] | wt5_sd_nan[41])}} & wt5_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[671:664] <= {8{(wt5_sd_nz[83] | wt5_sd_nan[41])}} & wt5_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[679:672] <= {8{(wt5_sd_nz[84] | wt5_sd_nan[42])}} & wt5_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[687:680] <= {8{(wt5_sd_nz[85] | wt5_sd_nan[42])}} & wt5_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[695:688] <= {8{(wt5_sd_nz[86] | wt5_sd_nan[43])}} & wt5_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[703:696] <= {8{(wt5_sd_nz[87] | wt5_sd_nan[43])}} & wt5_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[711:704] <= {8{(wt5_sd_nz[88] | wt5_sd_nan[44])}} & wt5_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[719:712] <= {8{(wt5_sd_nz[89] | wt5_sd_nan[44])}} & wt5_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[727:720] <= {8{(wt5_sd_nz[90] | wt5_sd_nan[45])}} & wt5_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[735:728] <= {8{(wt5_sd_nz[91] | wt5_sd_nan[45])}} & wt5_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[743:736] <= {8{(wt5_sd_nz[92] | wt5_sd_nan[46])}} & wt5_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[751:744] <= {8{(wt5_sd_nz[93] | wt5_sd_nan[46])}} & wt5_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[759:752] <= {8{(wt5_sd_nz[94] | wt5_sd_nan[47])}} & wt5_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[767:760] <= {8{(wt5_sd_nz[95] | wt5_sd_nan[47])}} & wt5_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[775:768] <= {8{(wt5_sd_nz[96] | wt5_sd_nan[48])}} & wt5_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[783:776] <= {8{(wt5_sd_nz[97] | wt5_sd_nan[48])}} & wt5_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[791:784] <= {8{(wt5_sd_nz[98] | wt5_sd_nan[49])}} & wt5_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[799:792] <= {8{(wt5_sd_nz[99] | wt5_sd_nan[49])}} & wt5_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[807:800] <= {8{(wt5_sd_nz[100] | wt5_sd_nan[50])}} & wt5_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[815:808] <= {8{(wt5_sd_nz[101] | wt5_sd_nan[50])}} & wt5_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[823:816] <= {8{(wt5_sd_nz[102] | wt5_sd_nan[51])}} & wt5_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[831:824] <= {8{(wt5_sd_nz[103] | wt5_sd_nan[51])}} & wt5_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[839:832] <= {8{(wt5_sd_nz[104] | wt5_sd_nan[52])}} & wt5_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[847:840] <= {8{(wt5_sd_nz[105] | wt5_sd_nan[52])}} & wt5_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[855:848] <= {8{(wt5_sd_nz[106] | wt5_sd_nan[53])}} & wt5_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[863:856] <= {8{(wt5_sd_nz[107] | wt5_sd_nan[53])}} & wt5_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[871:864] <= {8{(wt5_sd_nz[108] | wt5_sd_nan[54])}} & wt5_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[879:872] <= {8{(wt5_sd_nz[109] | wt5_sd_nan[54])}} & wt5_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[887:880] <= {8{(wt5_sd_nz[110] | wt5_sd_nan[55])}} & wt5_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[895:888] <= {8{(wt5_sd_nz[111] | wt5_sd_nan[55])}} & wt5_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[903:896] <= {8{(wt5_sd_nz[112] | wt5_sd_nan[56])}} & wt5_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[911:904] <= {8{(wt5_sd_nz[113] | wt5_sd_nan[56])}} & wt5_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[919:912] <= {8{(wt5_sd_nz[114] | wt5_sd_nan[57])}} & wt5_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[927:920] <= {8{(wt5_sd_nz[115] | wt5_sd_nan[57])}} & wt5_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[935:928] <= {8{(wt5_sd_nz[116] | wt5_sd_nan[58])}} & wt5_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[943:936] <= {8{(wt5_sd_nz[117] | wt5_sd_nan[58])}} & wt5_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[951:944] <= {8{(wt5_sd_nz[118] | wt5_sd_nan[59])}} & wt5_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[959:952] <= {8{(wt5_sd_nz[119] | wt5_sd_nan[59])}} & wt5_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[967:960] <= {8{(wt5_sd_nz[120] | wt5_sd_nan[60])}} & wt5_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[975:968] <= {8{(wt5_sd_nz[121] | wt5_sd_nan[60])}} & wt5_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[983:976] <= {8{(wt5_sd_nz[122] | wt5_sd_nan[61])}} & wt5_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[991:984] <= {8{(wt5_sd_nz[123] | wt5_sd_nan[61])}} & wt5_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[999:992] <= {8{(wt5_sd_nz[124] | wt5_sd_nan[62])}} & wt5_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[1007:1000] <= {8{(wt5_sd_nz[125] | wt5_sd_nan[62])}} & wt5_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[1015:1008] <= {8{(wt5_sd_nz[126] | wt5_sd_nan[63])}} & wt5_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b1) begin
    wt5_actv_data[1023:1016] <= {8{(wt5_sd_nz[127] | wt5_sd_nan[63])}} & wt5_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[5] & wt5_actv_pvld_w) == 1'b0) begin
  end else begin
    wt5_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt6_sd_pvld
  or dat_actv_stripe_end
  or wt6_actv_vld
  ) begin
    wt6_actv_pvld_w = dat_pre_stripe_st[6] ? wt6_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt6_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt6_actv_vld <= 1'b0;
  end else begin
  wt6_actv_vld <= wt6_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt6_actv_pvld <= {104{1'b0}};
  end else begin
  wt6_actv_pvld <= {104{wt6_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_nz <= wt6_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w & cfg_is_fp16_d1[80]) == 1'b1) begin
    wt6_actv_nan <= wt6_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w & cfg_is_fp16_d1[80]) == 1'b0) begin
  end else begin
    wt6_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[7:0] <= {8{(wt6_sd_nz[0] | wt6_sd_nan[0])}} & wt6_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[15:8] <= {8{(wt6_sd_nz[1] | wt6_sd_nan[0])}} & wt6_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[23:16] <= {8{(wt6_sd_nz[2] | wt6_sd_nan[1])}} & wt6_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[31:24] <= {8{(wt6_sd_nz[3] | wt6_sd_nan[1])}} & wt6_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[39:32] <= {8{(wt6_sd_nz[4] | wt6_sd_nan[2])}} & wt6_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[47:40] <= {8{(wt6_sd_nz[5] | wt6_sd_nan[2])}} & wt6_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[55:48] <= {8{(wt6_sd_nz[6] | wt6_sd_nan[3])}} & wt6_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[63:56] <= {8{(wt6_sd_nz[7] | wt6_sd_nan[3])}} & wt6_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[71:64] <= {8{(wt6_sd_nz[8] | wt6_sd_nan[4])}} & wt6_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[79:72] <= {8{(wt6_sd_nz[9] | wt6_sd_nan[4])}} & wt6_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[87:80] <= {8{(wt6_sd_nz[10] | wt6_sd_nan[5])}} & wt6_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[95:88] <= {8{(wt6_sd_nz[11] | wt6_sd_nan[5])}} & wt6_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[103:96] <= {8{(wt6_sd_nz[12] | wt6_sd_nan[6])}} & wt6_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[111:104] <= {8{(wt6_sd_nz[13] | wt6_sd_nan[6])}} & wt6_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[119:112] <= {8{(wt6_sd_nz[14] | wt6_sd_nan[7])}} & wt6_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[127:120] <= {8{(wt6_sd_nz[15] | wt6_sd_nan[7])}} & wt6_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[135:128] <= {8{(wt6_sd_nz[16] | wt6_sd_nan[8])}} & wt6_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[143:136] <= {8{(wt6_sd_nz[17] | wt6_sd_nan[8])}} & wt6_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[151:144] <= {8{(wt6_sd_nz[18] | wt6_sd_nan[9])}} & wt6_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[159:152] <= {8{(wt6_sd_nz[19] | wt6_sd_nan[9])}} & wt6_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[167:160] <= {8{(wt6_sd_nz[20] | wt6_sd_nan[10])}} & wt6_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[175:168] <= {8{(wt6_sd_nz[21] | wt6_sd_nan[10])}} & wt6_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[183:176] <= {8{(wt6_sd_nz[22] | wt6_sd_nan[11])}} & wt6_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[191:184] <= {8{(wt6_sd_nz[23] | wt6_sd_nan[11])}} & wt6_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[199:192] <= {8{(wt6_sd_nz[24] | wt6_sd_nan[12])}} & wt6_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[207:200] <= {8{(wt6_sd_nz[25] | wt6_sd_nan[12])}} & wt6_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[215:208] <= {8{(wt6_sd_nz[26] | wt6_sd_nan[13])}} & wt6_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[223:216] <= {8{(wt6_sd_nz[27] | wt6_sd_nan[13])}} & wt6_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[231:224] <= {8{(wt6_sd_nz[28] | wt6_sd_nan[14])}} & wt6_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[239:232] <= {8{(wt6_sd_nz[29] | wt6_sd_nan[14])}} & wt6_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[247:240] <= {8{(wt6_sd_nz[30] | wt6_sd_nan[15])}} & wt6_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[255:248] <= {8{(wt6_sd_nz[31] | wt6_sd_nan[15])}} & wt6_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[263:256] <= {8{(wt6_sd_nz[32] | wt6_sd_nan[16])}} & wt6_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[271:264] <= {8{(wt6_sd_nz[33] | wt6_sd_nan[16])}} & wt6_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[279:272] <= {8{(wt6_sd_nz[34] | wt6_sd_nan[17])}} & wt6_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[287:280] <= {8{(wt6_sd_nz[35] | wt6_sd_nan[17])}} & wt6_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[295:288] <= {8{(wt6_sd_nz[36] | wt6_sd_nan[18])}} & wt6_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[303:296] <= {8{(wt6_sd_nz[37] | wt6_sd_nan[18])}} & wt6_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[311:304] <= {8{(wt6_sd_nz[38] | wt6_sd_nan[19])}} & wt6_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[319:312] <= {8{(wt6_sd_nz[39] | wt6_sd_nan[19])}} & wt6_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[327:320] <= {8{(wt6_sd_nz[40] | wt6_sd_nan[20])}} & wt6_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[335:328] <= {8{(wt6_sd_nz[41] | wt6_sd_nan[20])}} & wt6_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[343:336] <= {8{(wt6_sd_nz[42] | wt6_sd_nan[21])}} & wt6_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[351:344] <= {8{(wt6_sd_nz[43] | wt6_sd_nan[21])}} & wt6_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[359:352] <= {8{(wt6_sd_nz[44] | wt6_sd_nan[22])}} & wt6_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[367:360] <= {8{(wt6_sd_nz[45] | wt6_sd_nan[22])}} & wt6_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[375:368] <= {8{(wt6_sd_nz[46] | wt6_sd_nan[23])}} & wt6_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[383:376] <= {8{(wt6_sd_nz[47] | wt6_sd_nan[23])}} & wt6_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[391:384] <= {8{(wt6_sd_nz[48] | wt6_sd_nan[24])}} & wt6_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[399:392] <= {8{(wt6_sd_nz[49] | wt6_sd_nan[24])}} & wt6_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[407:400] <= {8{(wt6_sd_nz[50] | wt6_sd_nan[25])}} & wt6_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[415:408] <= {8{(wt6_sd_nz[51] | wt6_sd_nan[25])}} & wt6_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[423:416] <= {8{(wt6_sd_nz[52] | wt6_sd_nan[26])}} & wt6_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[431:424] <= {8{(wt6_sd_nz[53] | wt6_sd_nan[26])}} & wt6_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[439:432] <= {8{(wt6_sd_nz[54] | wt6_sd_nan[27])}} & wt6_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[447:440] <= {8{(wt6_sd_nz[55] | wt6_sd_nan[27])}} & wt6_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[455:448] <= {8{(wt6_sd_nz[56] | wt6_sd_nan[28])}} & wt6_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[463:456] <= {8{(wt6_sd_nz[57] | wt6_sd_nan[28])}} & wt6_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[471:464] <= {8{(wt6_sd_nz[58] | wt6_sd_nan[29])}} & wt6_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[479:472] <= {8{(wt6_sd_nz[59] | wt6_sd_nan[29])}} & wt6_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[487:480] <= {8{(wt6_sd_nz[60] | wt6_sd_nan[30])}} & wt6_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[495:488] <= {8{(wt6_sd_nz[61] | wt6_sd_nan[30])}} & wt6_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[503:496] <= {8{(wt6_sd_nz[62] | wt6_sd_nan[31])}} & wt6_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[511:504] <= {8{(wt6_sd_nz[63] | wt6_sd_nan[31])}} & wt6_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[519:512] <= {8{(wt6_sd_nz[64] | wt6_sd_nan[32])}} & wt6_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[527:520] <= {8{(wt6_sd_nz[65] | wt6_sd_nan[32])}} & wt6_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[535:528] <= {8{(wt6_sd_nz[66] | wt6_sd_nan[33])}} & wt6_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[543:536] <= {8{(wt6_sd_nz[67] | wt6_sd_nan[33])}} & wt6_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[551:544] <= {8{(wt6_sd_nz[68] | wt6_sd_nan[34])}} & wt6_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[559:552] <= {8{(wt6_sd_nz[69] | wt6_sd_nan[34])}} & wt6_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[567:560] <= {8{(wt6_sd_nz[70] | wt6_sd_nan[35])}} & wt6_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[575:568] <= {8{(wt6_sd_nz[71] | wt6_sd_nan[35])}} & wt6_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[583:576] <= {8{(wt6_sd_nz[72] | wt6_sd_nan[36])}} & wt6_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[591:584] <= {8{(wt6_sd_nz[73] | wt6_sd_nan[36])}} & wt6_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[599:592] <= {8{(wt6_sd_nz[74] | wt6_sd_nan[37])}} & wt6_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[607:600] <= {8{(wt6_sd_nz[75] | wt6_sd_nan[37])}} & wt6_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[615:608] <= {8{(wt6_sd_nz[76] | wt6_sd_nan[38])}} & wt6_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[623:616] <= {8{(wt6_sd_nz[77] | wt6_sd_nan[38])}} & wt6_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[631:624] <= {8{(wt6_sd_nz[78] | wt6_sd_nan[39])}} & wt6_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[639:632] <= {8{(wt6_sd_nz[79] | wt6_sd_nan[39])}} & wt6_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[647:640] <= {8{(wt6_sd_nz[80] | wt6_sd_nan[40])}} & wt6_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[655:648] <= {8{(wt6_sd_nz[81] | wt6_sd_nan[40])}} & wt6_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[663:656] <= {8{(wt6_sd_nz[82] | wt6_sd_nan[41])}} & wt6_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[671:664] <= {8{(wt6_sd_nz[83] | wt6_sd_nan[41])}} & wt6_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[679:672] <= {8{(wt6_sd_nz[84] | wt6_sd_nan[42])}} & wt6_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[687:680] <= {8{(wt6_sd_nz[85] | wt6_sd_nan[42])}} & wt6_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[695:688] <= {8{(wt6_sd_nz[86] | wt6_sd_nan[43])}} & wt6_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[703:696] <= {8{(wt6_sd_nz[87] | wt6_sd_nan[43])}} & wt6_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[711:704] <= {8{(wt6_sd_nz[88] | wt6_sd_nan[44])}} & wt6_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[719:712] <= {8{(wt6_sd_nz[89] | wt6_sd_nan[44])}} & wt6_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[727:720] <= {8{(wt6_sd_nz[90] | wt6_sd_nan[45])}} & wt6_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[735:728] <= {8{(wt6_sd_nz[91] | wt6_sd_nan[45])}} & wt6_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[743:736] <= {8{(wt6_sd_nz[92] | wt6_sd_nan[46])}} & wt6_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[751:744] <= {8{(wt6_sd_nz[93] | wt6_sd_nan[46])}} & wt6_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[759:752] <= {8{(wt6_sd_nz[94] | wt6_sd_nan[47])}} & wt6_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[767:760] <= {8{(wt6_sd_nz[95] | wt6_sd_nan[47])}} & wt6_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[775:768] <= {8{(wt6_sd_nz[96] | wt6_sd_nan[48])}} & wt6_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[783:776] <= {8{(wt6_sd_nz[97] | wt6_sd_nan[48])}} & wt6_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[791:784] <= {8{(wt6_sd_nz[98] | wt6_sd_nan[49])}} & wt6_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[799:792] <= {8{(wt6_sd_nz[99] | wt6_sd_nan[49])}} & wt6_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[807:800] <= {8{(wt6_sd_nz[100] | wt6_sd_nan[50])}} & wt6_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[815:808] <= {8{(wt6_sd_nz[101] | wt6_sd_nan[50])}} & wt6_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[823:816] <= {8{(wt6_sd_nz[102] | wt6_sd_nan[51])}} & wt6_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[831:824] <= {8{(wt6_sd_nz[103] | wt6_sd_nan[51])}} & wt6_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[839:832] <= {8{(wt6_sd_nz[104] | wt6_sd_nan[52])}} & wt6_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[847:840] <= {8{(wt6_sd_nz[105] | wt6_sd_nan[52])}} & wt6_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[855:848] <= {8{(wt6_sd_nz[106] | wt6_sd_nan[53])}} & wt6_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[863:856] <= {8{(wt6_sd_nz[107] | wt6_sd_nan[53])}} & wt6_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[871:864] <= {8{(wt6_sd_nz[108] | wt6_sd_nan[54])}} & wt6_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[879:872] <= {8{(wt6_sd_nz[109] | wt6_sd_nan[54])}} & wt6_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[887:880] <= {8{(wt6_sd_nz[110] | wt6_sd_nan[55])}} & wt6_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[895:888] <= {8{(wt6_sd_nz[111] | wt6_sd_nan[55])}} & wt6_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[903:896] <= {8{(wt6_sd_nz[112] | wt6_sd_nan[56])}} & wt6_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[911:904] <= {8{(wt6_sd_nz[113] | wt6_sd_nan[56])}} & wt6_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[919:912] <= {8{(wt6_sd_nz[114] | wt6_sd_nan[57])}} & wt6_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[927:920] <= {8{(wt6_sd_nz[115] | wt6_sd_nan[57])}} & wt6_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[935:928] <= {8{(wt6_sd_nz[116] | wt6_sd_nan[58])}} & wt6_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[943:936] <= {8{(wt6_sd_nz[117] | wt6_sd_nan[58])}} & wt6_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[951:944] <= {8{(wt6_sd_nz[118] | wt6_sd_nan[59])}} & wt6_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[959:952] <= {8{(wt6_sd_nz[119] | wt6_sd_nan[59])}} & wt6_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[967:960] <= {8{(wt6_sd_nz[120] | wt6_sd_nan[60])}} & wt6_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[975:968] <= {8{(wt6_sd_nz[121] | wt6_sd_nan[60])}} & wt6_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[983:976] <= {8{(wt6_sd_nz[122] | wt6_sd_nan[61])}} & wt6_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[991:984] <= {8{(wt6_sd_nz[123] | wt6_sd_nan[61])}} & wt6_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[999:992] <= {8{(wt6_sd_nz[124] | wt6_sd_nan[62])}} & wt6_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[1007:1000] <= {8{(wt6_sd_nz[125] | wt6_sd_nan[62])}} & wt6_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[1015:1008] <= {8{(wt6_sd_nz[126] | wt6_sd_nan[63])}} & wt6_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b1) begin
    wt6_actv_data[1023:1016] <= {8{(wt6_sd_nz[127] | wt6_sd_nan[63])}} & wt6_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[6] & wt6_actv_pvld_w) == 1'b0) begin
  end else begin
    wt6_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(
  dat_pre_stripe_st
  or wt7_sd_pvld
  or dat_actv_stripe_end
  or wt7_actv_vld
  ) begin
    wt7_actv_pvld_w = dat_pre_stripe_st[7] ? wt7_sd_pvld :
                      dat_actv_stripe_end ? 1'b0 :
                      wt7_actv_vld[0];
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt7_actv_vld <= 1'b0;
  end else begin
  wt7_actv_vld <= wt7_actv_pvld_w;
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    wt7_actv_pvld <= {104{1'b0}};
  end else begin
  wt7_actv_pvld <= {104{wt7_actv_pvld_w}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_nz <= wt7_sd_nz;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w & cfg_is_fp16_d1[81]) == 1'b1) begin
    wt7_actv_nan <= wt7_sd_nan;
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w & cfg_is_fp16_d1[81]) == 1'b0) begin
  end else begin
    wt7_actv_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[7:0] <= {8{(wt7_sd_nz[0] | wt7_sd_nan[0])}} & wt7_sd_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[15:8] <= {8{(wt7_sd_nz[1] | wt7_sd_nan[0])}} & wt7_sd_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[23:16] <= {8{(wt7_sd_nz[2] | wt7_sd_nan[1])}} & wt7_sd_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[31:24] <= {8{(wt7_sd_nz[3] | wt7_sd_nan[1])}} & wt7_sd_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[39:32] <= {8{(wt7_sd_nz[4] | wt7_sd_nan[2])}} & wt7_sd_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[47:40] <= {8{(wt7_sd_nz[5] | wt7_sd_nan[2])}} & wt7_sd_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[55:48] <= {8{(wt7_sd_nz[6] | wt7_sd_nan[3])}} & wt7_sd_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[63:56] <= {8{(wt7_sd_nz[7] | wt7_sd_nan[3])}} & wt7_sd_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[71:64] <= {8{(wt7_sd_nz[8] | wt7_sd_nan[4])}} & wt7_sd_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[79:72] <= {8{(wt7_sd_nz[9] | wt7_sd_nan[4])}} & wt7_sd_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[87:80] <= {8{(wt7_sd_nz[10] | wt7_sd_nan[5])}} & wt7_sd_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[95:88] <= {8{(wt7_sd_nz[11] | wt7_sd_nan[5])}} & wt7_sd_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[103:96] <= {8{(wt7_sd_nz[12] | wt7_sd_nan[6])}} & wt7_sd_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[111:104] <= {8{(wt7_sd_nz[13] | wt7_sd_nan[6])}} & wt7_sd_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[119:112] <= {8{(wt7_sd_nz[14] | wt7_sd_nan[7])}} & wt7_sd_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[127:120] <= {8{(wt7_sd_nz[15] | wt7_sd_nan[7])}} & wt7_sd_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[135:128] <= {8{(wt7_sd_nz[16] | wt7_sd_nan[8])}} & wt7_sd_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[143:136] <= {8{(wt7_sd_nz[17] | wt7_sd_nan[8])}} & wt7_sd_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[151:144] <= {8{(wt7_sd_nz[18] | wt7_sd_nan[9])}} & wt7_sd_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[159:152] <= {8{(wt7_sd_nz[19] | wt7_sd_nan[9])}} & wt7_sd_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[167:160] <= {8{(wt7_sd_nz[20] | wt7_sd_nan[10])}} & wt7_sd_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[175:168] <= {8{(wt7_sd_nz[21] | wt7_sd_nan[10])}} & wt7_sd_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[183:176] <= {8{(wt7_sd_nz[22] | wt7_sd_nan[11])}} & wt7_sd_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[191:184] <= {8{(wt7_sd_nz[23] | wt7_sd_nan[11])}} & wt7_sd_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[199:192] <= {8{(wt7_sd_nz[24] | wt7_sd_nan[12])}} & wt7_sd_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[207:200] <= {8{(wt7_sd_nz[25] | wt7_sd_nan[12])}} & wt7_sd_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[215:208] <= {8{(wt7_sd_nz[26] | wt7_sd_nan[13])}} & wt7_sd_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[223:216] <= {8{(wt7_sd_nz[27] | wt7_sd_nan[13])}} & wt7_sd_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[231:224] <= {8{(wt7_sd_nz[28] | wt7_sd_nan[14])}} & wt7_sd_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[239:232] <= {8{(wt7_sd_nz[29] | wt7_sd_nan[14])}} & wt7_sd_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[247:240] <= {8{(wt7_sd_nz[30] | wt7_sd_nan[15])}} & wt7_sd_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[255:248] <= {8{(wt7_sd_nz[31] | wt7_sd_nan[15])}} & wt7_sd_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[263:256] <= {8{(wt7_sd_nz[32] | wt7_sd_nan[16])}} & wt7_sd_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[271:264] <= {8{(wt7_sd_nz[33] | wt7_sd_nan[16])}} & wt7_sd_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[279:272] <= {8{(wt7_sd_nz[34] | wt7_sd_nan[17])}} & wt7_sd_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[287:280] <= {8{(wt7_sd_nz[35] | wt7_sd_nan[17])}} & wt7_sd_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[295:288] <= {8{(wt7_sd_nz[36] | wt7_sd_nan[18])}} & wt7_sd_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[303:296] <= {8{(wt7_sd_nz[37] | wt7_sd_nan[18])}} & wt7_sd_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[311:304] <= {8{(wt7_sd_nz[38] | wt7_sd_nan[19])}} & wt7_sd_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[319:312] <= {8{(wt7_sd_nz[39] | wt7_sd_nan[19])}} & wt7_sd_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[327:320] <= {8{(wt7_sd_nz[40] | wt7_sd_nan[20])}} & wt7_sd_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[335:328] <= {8{(wt7_sd_nz[41] | wt7_sd_nan[20])}} & wt7_sd_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[343:336] <= {8{(wt7_sd_nz[42] | wt7_sd_nan[21])}} & wt7_sd_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[351:344] <= {8{(wt7_sd_nz[43] | wt7_sd_nan[21])}} & wt7_sd_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[359:352] <= {8{(wt7_sd_nz[44] | wt7_sd_nan[22])}} & wt7_sd_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[367:360] <= {8{(wt7_sd_nz[45] | wt7_sd_nan[22])}} & wt7_sd_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[375:368] <= {8{(wt7_sd_nz[46] | wt7_sd_nan[23])}} & wt7_sd_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[383:376] <= {8{(wt7_sd_nz[47] | wt7_sd_nan[23])}} & wt7_sd_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[391:384] <= {8{(wt7_sd_nz[48] | wt7_sd_nan[24])}} & wt7_sd_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[399:392] <= {8{(wt7_sd_nz[49] | wt7_sd_nan[24])}} & wt7_sd_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[407:400] <= {8{(wt7_sd_nz[50] | wt7_sd_nan[25])}} & wt7_sd_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[415:408] <= {8{(wt7_sd_nz[51] | wt7_sd_nan[25])}} & wt7_sd_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[423:416] <= {8{(wt7_sd_nz[52] | wt7_sd_nan[26])}} & wt7_sd_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[431:424] <= {8{(wt7_sd_nz[53] | wt7_sd_nan[26])}} & wt7_sd_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[439:432] <= {8{(wt7_sd_nz[54] | wt7_sd_nan[27])}} & wt7_sd_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[447:440] <= {8{(wt7_sd_nz[55] | wt7_sd_nan[27])}} & wt7_sd_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[455:448] <= {8{(wt7_sd_nz[56] | wt7_sd_nan[28])}} & wt7_sd_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[463:456] <= {8{(wt7_sd_nz[57] | wt7_sd_nan[28])}} & wt7_sd_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[471:464] <= {8{(wt7_sd_nz[58] | wt7_sd_nan[29])}} & wt7_sd_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[479:472] <= {8{(wt7_sd_nz[59] | wt7_sd_nan[29])}} & wt7_sd_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[487:480] <= {8{(wt7_sd_nz[60] | wt7_sd_nan[30])}} & wt7_sd_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[495:488] <= {8{(wt7_sd_nz[61] | wt7_sd_nan[30])}} & wt7_sd_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[503:496] <= {8{(wt7_sd_nz[62] | wt7_sd_nan[31])}} & wt7_sd_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[511:504] <= {8{(wt7_sd_nz[63] | wt7_sd_nan[31])}} & wt7_sd_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[519:512] <= {8{(wt7_sd_nz[64] | wt7_sd_nan[32])}} & wt7_sd_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[527:520] <= {8{(wt7_sd_nz[65] | wt7_sd_nan[32])}} & wt7_sd_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[535:528] <= {8{(wt7_sd_nz[66] | wt7_sd_nan[33])}} & wt7_sd_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[543:536] <= {8{(wt7_sd_nz[67] | wt7_sd_nan[33])}} & wt7_sd_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[551:544] <= {8{(wt7_sd_nz[68] | wt7_sd_nan[34])}} & wt7_sd_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[559:552] <= {8{(wt7_sd_nz[69] | wt7_sd_nan[34])}} & wt7_sd_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[567:560] <= {8{(wt7_sd_nz[70] | wt7_sd_nan[35])}} & wt7_sd_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[575:568] <= {8{(wt7_sd_nz[71] | wt7_sd_nan[35])}} & wt7_sd_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[583:576] <= {8{(wt7_sd_nz[72] | wt7_sd_nan[36])}} & wt7_sd_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[591:584] <= {8{(wt7_sd_nz[73] | wt7_sd_nan[36])}} & wt7_sd_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[599:592] <= {8{(wt7_sd_nz[74] | wt7_sd_nan[37])}} & wt7_sd_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[607:600] <= {8{(wt7_sd_nz[75] | wt7_sd_nan[37])}} & wt7_sd_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[615:608] <= {8{(wt7_sd_nz[76] | wt7_sd_nan[38])}} & wt7_sd_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[623:616] <= {8{(wt7_sd_nz[77] | wt7_sd_nan[38])}} & wt7_sd_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[631:624] <= {8{(wt7_sd_nz[78] | wt7_sd_nan[39])}} & wt7_sd_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[639:632] <= {8{(wt7_sd_nz[79] | wt7_sd_nan[39])}} & wt7_sd_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[647:640] <= {8{(wt7_sd_nz[80] | wt7_sd_nan[40])}} & wt7_sd_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[655:648] <= {8{(wt7_sd_nz[81] | wt7_sd_nan[40])}} & wt7_sd_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[663:656] <= {8{(wt7_sd_nz[82] | wt7_sd_nan[41])}} & wt7_sd_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[671:664] <= {8{(wt7_sd_nz[83] | wt7_sd_nan[41])}} & wt7_sd_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[679:672] <= {8{(wt7_sd_nz[84] | wt7_sd_nan[42])}} & wt7_sd_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[687:680] <= {8{(wt7_sd_nz[85] | wt7_sd_nan[42])}} & wt7_sd_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[695:688] <= {8{(wt7_sd_nz[86] | wt7_sd_nan[43])}} & wt7_sd_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[703:696] <= {8{(wt7_sd_nz[87] | wt7_sd_nan[43])}} & wt7_sd_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[711:704] <= {8{(wt7_sd_nz[88] | wt7_sd_nan[44])}} & wt7_sd_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[719:712] <= {8{(wt7_sd_nz[89] | wt7_sd_nan[44])}} & wt7_sd_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[727:720] <= {8{(wt7_sd_nz[90] | wt7_sd_nan[45])}} & wt7_sd_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[735:728] <= {8{(wt7_sd_nz[91] | wt7_sd_nan[45])}} & wt7_sd_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[743:736] <= {8{(wt7_sd_nz[92] | wt7_sd_nan[46])}} & wt7_sd_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[751:744] <= {8{(wt7_sd_nz[93] | wt7_sd_nan[46])}} & wt7_sd_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[759:752] <= {8{(wt7_sd_nz[94] | wt7_sd_nan[47])}} & wt7_sd_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[767:760] <= {8{(wt7_sd_nz[95] | wt7_sd_nan[47])}} & wt7_sd_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[775:768] <= {8{(wt7_sd_nz[96] | wt7_sd_nan[48])}} & wt7_sd_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[783:776] <= {8{(wt7_sd_nz[97] | wt7_sd_nan[48])}} & wt7_sd_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[791:784] <= {8{(wt7_sd_nz[98] | wt7_sd_nan[49])}} & wt7_sd_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[799:792] <= {8{(wt7_sd_nz[99] | wt7_sd_nan[49])}} & wt7_sd_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[807:800] <= {8{(wt7_sd_nz[100] | wt7_sd_nan[50])}} & wt7_sd_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[815:808] <= {8{(wt7_sd_nz[101] | wt7_sd_nan[50])}} & wt7_sd_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[823:816] <= {8{(wt7_sd_nz[102] | wt7_sd_nan[51])}} & wt7_sd_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[831:824] <= {8{(wt7_sd_nz[103] | wt7_sd_nan[51])}} & wt7_sd_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[839:832] <= {8{(wt7_sd_nz[104] | wt7_sd_nan[52])}} & wt7_sd_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[847:840] <= {8{(wt7_sd_nz[105] | wt7_sd_nan[52])}} & wt7_sd_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[855:848] <= {8{(wt7_sd_nz[106] | wt7_sd_nan[53])}} & wt7_sd_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[863:856] <= {8{(wt7_sd_nz[107] | wt7_sd_nan[53])}} & wt7_sd_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[871:864] <= {8{(wt7_sd_nz[108] | wt7_sd_nan[54])}} & wt7_sd_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[879:872] <= {8{(wt7_sd_nz[109] | wt7_sd_nan[54])}} & wt7_sd_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[887:880] <= {8{(wt7_sd_nz[110] | wt7_sd_nan[55])}} & wt7_sd_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[895:888] <= {8{(wt7_sd_nz[111] | wt7_sd_nan[55])}} & wt7_sd_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[903:896] <= {8{(wt7_sd_nz[112] | wt7_sd_nan[56])}} & wt7_sd_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[911:904] <= {8{(wt7_sd_nz[113] | wt7_sd_nan[56])}} & wt7_sd_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[919:912] <= {8{(wt7_sd_nz[114] | wt7_sd_nan[57])}} & wt7_sd_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[927:920] <= {8{(wt7_sd_nz[115] | wt7_sd_nan[57])}} & wt7_sd_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[935:928] <= {8{(wt7_sd_nz[116] | wt7_sd_nan[58])}} & wt7_sd_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[943:936] <= {8{(wt7_sd_nz[117] | wt7_sd_nan[58])}} & wt7_sd_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[951:944] <= {8{(wt7_sd_nz[118] | wt7_sd_nan[59])}} & wt7_sd_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[959:952] <= {8{(wt7_sd_nz[119] | wt7_sd_nan[59])}} & wt7_sd_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[967:960] <= {8{(wt7_sd_nz[120] | wt7_sd_nan[60])}} & wt7_sd_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[975:968] <= {8{(wt7_sd_nz[121] | wt7_sd_nan[60])}} & wt7_sd_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[983:976] <= {8{(wt7_sd_nz[122] | wt7_sd_nan[61])}} & wt7_sd_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[991:984] <= {8{(wt7_sd_nz[123] | wt7_sd_nan[61])}} & wt7_sd_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[999:992] <= {8{(wt7_sd_nz[124] | wt7_sd_nan[62])}} & wt7_sd_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[1007:1000] <= {8{(wt7_sd_nz[125] | wt7_sd_nan[62])}} & wt7_sd_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[1015:1008] <= {8{(wt7_sd_nz[126] | wt7_sd_nan[63])}} & wt7_sd_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b1) begin
    wt7_actv_data[1023:1016] <= {8{(wt7_sd_nz[127] | wt7_sd_nan[63])}} & wt7_sd_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_stripe_st[7] & wt7_actv_pvld_w) == 1'b0) begin
  end else begin
    wt7_actv_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt0_active_pvld conflict!")      zzz_assert_never_4x (nvdla_core_clk, `ASSERT_RESET, (wt0_sd_pvld & wt_pre_sel[0] & ~dat_pre_stripe_st[0])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt1_active_pvld conflict!")      zzz_assert_never_5x (nvdla_core_clk, `ASSERT_RESET, (wt1_sd_pvld & wt_pre_sel[1] & ~dat_pre_stripe_st[1])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt2_active_pvld conflict!")      zzz_assert_never_6x (nvdla_core_clk, `ASSERT_RESET, (wt2_sd_pvld & wt_pre_sel[2] & ~dat_pre_stripe_st[2])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt3_active_pvld conflict!")      zzz_assert_never_7x (nvdla_core_clk, `ASSERT_RESET, (wt3_sd_pvld & wt_pre_sel[3] & ~dat_pre_stripe_st[3])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt4_active_pvld conflict!")      zzz_assert_never_8x (nvdla_core_clk, `ASSERT_RESET, (wt4_sd_pvld & wt_pre_sel[4] & ~dat_pre_stripe_st[4])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt5_active_pvld conflict!")      zzz_assert_never_9x (nvdla_core_clk, `ASSERT_RESET, (wt5_sd_pvld & wt_pre_sel[5] & ~dat_pre_stripe_st[5])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt6_active_pvld conflict!")      zzz_assert_never_10x (nvdla_core_clk, `ASSERT_RESET, (wt6_sd_pvld & wt_pre_sel[6] & ~dat_pre_stripe_st[6])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML 
// spyglass disable_block STARC-2.10.3.2a 
// spyglass disable_block STARC05-2.1.3.1 
// spyglass disable_block STARC-2.1.4.6 
// spyglass disable_block W116 
// spyglass disable_block W154 
// spyglass disable_block W239 
// spyglass disable_block W362 
// spyglass disable_block WRN_58 
// spyglass disable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET nvdla_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b0 : nvdla_core_rstn)
`else
`define ASSERT_RESET ((1'bx === nvdla_core_rstn) ? 1'b1 : nvdla_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
  // VCS coverage off 
  nv_assert_never #(0,0,"Error! wt7_active_pvld conflict!")      zzz_assert_never_11x (nvdla_core_clk, `ASSERT_RESET, (wt7_sd_pvld & wt_pre_sel[7] & ~dat_pre_stripe_st[7])); // spyglass disable W504 SelfDeterminedExpr-ML 
  // VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML 
// spyglass enable_block STARC-2.10.3.2a 
// spyglass enable_block STARC05-2.1.3.1 
// spyglass enable_block STARC-2.1.4.6 
// spyglass enable_block W116 
// spyglass enable_block W154 
// spyglass enable_block W239 
// spyglass enable_block W362 
// spyglass enable_block WRN_58 
// spyglass enable_block WRN_61 
`endif // SPYGLASS_ASSERT_ON



always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_stripe_end <= 1'b0;
  end else begin
  dat_actv_stripe_end <= dat_pre_stripe_end[8];
  end
end

//==========================================================
// Data reordering and detect
//==========================================================

always @(
  in_dat_data127
  or in_dat_data126
  or in_dat_data125
  or in_dat_data124
  or in_dat_data123
  or in_dat_data122
  or in_dat_data121
  or in_dat_data120
  or in_dat_data119
  or in_dat_data118
  or in_dat_data117
  or in_dat_data116
  or in_dat_data115
  or in_dat_data114
  or in_dat_data113
  or in_dat_data112
  or in_dat_data111
  or in_dat_data110
  or in_dat_data109
  or in_dat_data108
  or in_dat_data107
  or in_dat_data106
  or in_dat_data105
  or in_dat_data104
  or in_dat_data103
  or in_dat_data102
  or in_dat_data101
  or in_dat_data100
  or in_dat_data99
  or in_dat_data98
  or in_dat_data97
  or in_dat_data96
  or in_dat_data95
  or in_dat_data94
  or in_dat_data93
  or in_dat_data92
  or in_dat_data91
  or in_dat_data90
  or in_dat_data89
  or in_dat_data88
  or in_dat_data87
  or in_dat_data86
  or in_dat_data85
  or in_dat_data84
  or in_dat_data83
  or in_dat_data82
  or in_dat_data81
  or in_dat_data80
  or in_dat_data79
  or in_dat_data78
  or in_dat_data77
  or in_dat_data76
  or in_dat_data75
  or in_dat_data74
  or in_dat_data73
  or in_dat_data72
  or in_dat_data71
  or in_dat_data70
  or in_dat_data69
  or in_dat_data68
  or in_dat_data67
  or in_dat_data66
  or in_dat_data65
  or in_dat_data64
  or in_dat_data63
  or in_dat_data62
  or in_dat_data61
  or in_dat_data60
  or in_dat_data59
  or in_dat_data58
  or in_dat_data57
  or in_dat_data56
  or in_dat_data55
  or in_dat_data54
  or in_dat_data53
  or in_dat_data52
  or in_dat_data51
  or in_dat_data50
  or in_dat_data49
  or in_dat_data48
  or in_dat_data47
  or in_dat_data46
  or in_dat_data45
  or in_dat_data44
  or in_dat_data43
  or in_dat_data42
  or in_dat_data41
  or in_dat_data40
  or in_dat_data39
  or in_dat_data38
  or in_dat_data37
  or in_dat_data36
  or in_dat_data35
  or in_dat_data34
  or in_dat_data33
  or in_dat_data32
  or in_dat_data31
  or in_dat_data30
  or in_dat_data29
  or in_dat_data28
  or in_dat_data27
  or in_dat_data26
  or in_dat_data25
  or in_dat_data24
  or in_dat_data23
  or in_dat_data22
  or in_dat_data21
  or in_dat_data20
  or in_dat_data19
  or in_dat_data18
  or in_dat_data17
  or in_dat_data16
  or in_dat_data15
  or in_dat_data14
  or in_dat_data13
  or in_dat_data12
  or in_dat_data11
  or in_dat_data10
  or in_dat_data9
  or in_dat_data8
  or in_dat_data7
  or in_dat_data6
  or in_dat_data5
  or in_dat_data4
  or in_dat_data3
  or in_dat_data2
  or in_dat_data1
  or in_dat_data0
  ) begin
    in_dat_data_pack = {in_dat_data127, in_dat_data126, in_dat_data125, in_dat_data124, in_dat_data123, in_dat_data122, in_dat_data121, in_dat_data120, in_dat_data119, in_dat_data118, in_dat_data117, in_dat_data116, in_dat_data115, in_dat_data114, in_dat_data113, in_dat_data112, in_dat_data111, in_dat_data110, in_dat_data109, in_dat_data108, in_dat_data107, in_dat_data106, in_dat_data105, in_dat_data104, in_dat_data103, in_dat_data102, in_dat_data101, in_dat_data100, in_dat_data99, in_dat_data98, in_dat_data97, in_dat_data96, in_dat_data95, in_dat_data94, in_dat_data93, in_dat_data92, in_dat_data91, in_dat_data90, in_dat_data89, in_dat_data88, in_dat_data87, in_dat_data86, in_dat_data85, in_dat_data84, in_dat_data83, in_dat_data82, in_dat_data81, in_dat_data80, in_dat_data79, in_dat_data78, in_dat_data77, in_dat_data76, in_dat_data75, in_dat_data74, in_dat_data73, in_dat_data72, in_dat_data71, in_dat_data70, in_dat_data69, in_dat_data68, in_dat_data67, in_dat_data66, in_dat_data65, in_dat_data64, in_dat_data63, in_dat_data62, in_dat_data61, in_dat_data60, in_dat_data59, in_dat_data58, in_dat_data57, in_dat_data56, in_dat_data55, in_dat_data54, in_dat_data53, in_dat_data52, in_dat_data51, in_dat_data50, in_dat_data49, in_dat_data48, in_dat_data47, in_dat_data46, in_dat_data45, in_dat_data44, in_dat_data43, in_dat_data42, in_dat_data41, in_dat_data40, in_dat_data39, in_dat_data38, in_dat_data37, in_dat_data36, in_dat_data35, in_dat_data34, in_dat_data33, in_dat_data32, in_dat_data31, in_dat_data30, in_dat_data29, in_dat_data28, in_dat_data27, in_dat_data26, in_dat_data25, in_dat_data24, in_dat_data23, in_dat_data22, in_dat_data21, in_dat_data20, in_dat_data19, in_dat_data18, in_dat_data17, in_dat_data16, in_dat_data15, in_dat_data14, in_dat_data13, in_dat_data12, in_dat_data11, in_dat_data10, in_dat_data9, in_dat_data8, in_dat_data7, in_dat_data6, in_dat_data5, in_dat_data4, in_dat_data3, in_dat_data2, in_dat_data1, in_dat_data0};
end

//////////////// in_wt_data_int16 ////////////////
always @(
  cfg_is_int16_d1
  or in_dat_data127
  or in_dat_data126
  or in_dat_data125
  or in_dat_data124
  or in_dat_data123
  or in_dat_data122
  or in_dat_data121
  or in_dat_data120
  or in_dat_data119
  or in_dat_data118
  or in_dat_data117
  or in_dat_data116
  or in_dat_data115
  or in_dat_data114
  or in_dat_data113
  or in_dat_data112
  or in_dat_data111
  or in_dat_data110
  or in_dat_data109
  or in_dat_data108
  or in_dat_data107
  or in_dat_data106
  or in_dat_data105
  or in_dat_data104
  or in_dat_data103
  or in_dat_data102
  or in_dat_data101
  or in_dat_data100
  or in_dat_data99
  or in_dat_data98
  or in_dat_data97
  or in_dat_data96
  or in_dat_data95
  or in_dat_data94
  or in_dat_data93
  or in_dat_data92
  or in_dat_data91
  or in_dat_data90
  or in_dat_data89
  or in_dat_data88
  or in_dat_data87
  or in_dat_data86
  or in_dat_data85
  or in_dat_data84
  or in_dat_data83
  or in_dat_data82
  or in_dat_data81
  or in_dat_data80
  or in_dat_data79
  or in_dat_data78
  or in_dat_data77
  or in_dat_data76
  or in_dat_data75
  or in_dat_data74
  or in_dat_data73
  or in_dat_data72
  or in_dat_data71
  or in_dat_data70
  or in_dat_data69
  or in_dat_data68
  or in_dat_data67
  or in_dat_data66
  or in_dat_data65
  or in_dat_data64
  or in_dat_data63
  or in_dat_data62
  or in_dat_data61
  or in_dat_data60
  or in_dat_data59
  or in_dat_data58
  or in_dat_data57
  or in_dat_data56
  or in_dat_data55
  or in_dat_data54
  or in_dat_data53
  or in_dat_data52
  or in_dat_data51
  or in_dat_data50
  or in_dat_data49
  or in_dat_data48
  or in_dat_data47
  or in_dat_data46
  or in_dat_data45
  or in_dat_data44
  or in_dat_data43
  or in_dat_data42
  or in_dat_data41
  or in_dat_data40
  or in_dat_data39
  or in_dat_data38
  or in_dat_data37
  or in_dat_data36
  or in_dat_data35
  or in_dat_data34
  or in_dat_data33
  or in_dat_data32
  or in_dat_data31
  or in_dat_data30
  or in_dat_data29
  or in_dat_data28
  or in_dat_data27
  or in_dat_data26
  or in_dat_data25
  or in_dat_data24
  or in_dat_data23
  or in_dat_data22
  or in_dat_data21
  or in_dat_data20
  or in_dat_data19
  or in_dat_data18
  or in_dat_data17
  or in_dat_data16
  or in_dat_data15
  or in_dat_data14
  or in_dat_data13
  or in_dat_data12
  or in_dat_data11
  or in_dat_data10
  or in_dat_data9
  or in_dat_data8
  or in_dat_data7
  or in_dat_data6
  or in_dat_data5
  or in_dat_data4
  or in_dat_data3
  or in_dat_data2
  or in_dat_data1
  or in_dat_data0
  ) begin
    in_dat_data_int16_63 = ({16{cfg_is_int16_d1[63]}} & {in_dat_data127, in_dat_data126});
    in_dat_data_int16_62 = ({16{cfg_is_int16_d1[62]}} & {in_dat_data125, in_dat_data124});
    in_dat_data_int16_61 = ({16{cfg_is_int16_d1[61]}} & {in_dat_data123, in_dat_data122});
    in_dat_data_int16_60 = ({16{cfg_is_int16_d1[60]}} & {in_dat_data121, in_dat_data120});
    in_dat_data_int16_59 = ({16{cfg_is_int16_d1[59]}} & {in_dat_data119, in_dat_data118});
    in_dat_data_int16_58 = ({16{cfg_is_int16_d1[58]}} & {in_dat_data117, in_dat_data116});
    in_dat_data_int16_57 = ({16{cfg_is_int16_d1[57]}} & {in_dat_data115, in_dat_data114});
    in_dat_data_int16_56 = ({16{cfg_is_int16_d1[56]}} & {in_dat_data113, in_dat_data112});
    in_dat_data_int16_55 = ({16{cfg_is_int16_d1[55]}} & {in_dat_data111, in_dat_data110});
    in_dat_data_int16_54 = ({16{cfg_is_int16_d1[54]}} & {in_dat_data109, in_dat_data108});
    in_dat_data_int16_53 = ({16{cfg_is_int16_d1[53]}} & {in_dat_data107, in_dat_data106});
    in_dat_data_int16_52 = ({16{cfg_is_int16_d1[52]}} & {in_dat_data105, in_dat_data104});
    in_dat_data_int16_51 = ({16{cfg_is_int16_d1[51]}} & {in_dat_data103, in_dat_data102});
    in_dat_data_int16_50 = ({16{cfg_is_int16_d1[50]}} & {in_dat_data101, in_dat_data100});
    in_dat_data_int16_49 = ({16{cfg_is_int16_d1[49]}} & {in_dat_data99, in_dat_data98});
    in_dat_data_int16_48 = ({16{cfg_is_int16_d1[48]}} & {in_dat_data97, in_dat_data96});
    in_dat_data_int16_47 = ({16{cfg_is_int16_d1[47]}} & {in_dat_data95, in_dat_data94});
    in_dat_data_int16_46 = ({16{cfg_is_int16_d1[46]}} & {in_dat_data93, in_dat_data92});
    in_dat_data_int16_45 = ({16{cfg_is_int16_d1[45]}} & {in_dat_data91, in_dat_data90});
    in_dat_data_int16_44 = ({16{cfg_is_int16_d1[44]}} & {in_dat_data89, in_dat_data88});
    in_dat_data_int16_43 = ({16{cfg_is_int16_d1[43]}} & {in_dat_data87, in_dat_data86});
    in_dat_data_int16_42 = ({16{cfg_is_int16_d1[42]}} & {in_dat_data85, in_dat_data84});
    in_dat_data_int16_41 = ({16{cfg_is_int16_d1[41]}} & {in_dat_data83, in_dat_data82});
    in_dat_data_int16_40 = ({16{cfg_is_int16_d1[40]}} & {in_dat_data81, in_dat_data80});
    in_dat_data_int16_39 = ({16{cfg_is_int16_d1[39]}} & {in_dat_data79, in_dat_data78});
    in_dat_data_int16_38 = ({16{cfg_is_int16_d1[38]}} & {in_dat_data77, in_dat_data76});
    in_dat_data_int16_37 = ({16{cfg_is_int16_d1[37]}} & {in_dat_data75, in_dat_data74});
    in_dat_data_int16_36 = ({16{cfg_is_int16_d1[36]}} & {in_dat_data73, in_dat_data72});
    in_dat_data_int16_35 = ({16{cfg_is_int16_d1[35]}} & {in_dat_data71, in_dat_data70});
    in_dat_data_int16_34 = ({16{cfg_is_int16_d1[34]}} & {in_dat_data69, in_dat_data68});
    in_dat_data_int16_33 = ({16{cfg_is_int16_d1[33]}} & {in_dat_data67, in_dat_data66});
    in_dat_data_int16_32 = ({16{cfg_is_int16_d1[32]}} & {in_dat_data65, in_dat_data64});
    in_dat_data_int16_31 = ({16{cfg_is_int16_d1[31]}} & {in_dat_data63, in_dat_data62});
    in_dat_data_int16_30 = ({16{cfg_is_int16_d1[30]}} & {in_dat_data61, in_dat_data60});
    in_dat_data_int16_29 = ({16{cfg_is_int16_d1[29]}} & {in_dat_data59, in_dat_data58});
    in_dat_data_int16_28 = ({16{cfg_is_int16_d1[28]}} & {in_dat_data57, in_dat_data56});
    in_dat_data_int16_27 = ({16{cfg_is_int16_d1[27]}} & {in_dat_data55, in_dat_data54});
    in_dat_data_int16_26 = ({16{cfg_is_int16_d1[26]}} & {in_dat_data53, in_dat_data52});
    in_dat_data_int16_25 = ({16{cfg_is_int16_d1[25]}} & {in_dat_data51, in_dat_data50});
    in_dat_data_int16_24 = ({16{cfg_is_int16_d1[24]}} & {in_dat_data49, in_dat_data48});
    in_dat_data_int16_23 = ({16{cfg_is_int16_d1[23]}} & {in_dat_data47, in_dat_data46});
    in_dat_data_int16_22 = ({16{cfg_is_int16_d1[22]}} & {in_dat_data45, in_dat_data44});
    in_dat_data_int16_21 = ({16{cfg_is_int16_d1[21]}} & {in_dat_data43, in_dat_data42});
    in_dat_data_int16_20 = ({16{cfg_is_int16_d1[20]}} & {in_dat_data41, in_dat_data40});
    in_dat_data_int16_19 = ({16{cfg_is_int16_d1[19]}} & {in_dat_data39, in_dat_data38});
    in_dat_data_int16_18 = ({16{cfg_is_int16_d1[18]}} & {in_dat_data37, in_dat_data36});
    in_dat_data_int16_17 = ({16{cfg_is_int16_d1[17]}} & {in_dat_data35, in_dat_data34});
    in_dat_data_int16_16 = ({16{cfg_is_int16_d1[16]}} & {in_dat_data33, in_dat_data32});
    in_dat_data_int16_15 = ({16{cfg_is_int16_d1[15]}} & {in_dat_data31, in_dat_data30});
    in_dat_data_int16_14 = ({16{cfg_is_int16_d1[14]}} & {in_dat_data29, in_dat_data28});
    in_dat_data_int16_13 = ({16{cfg_is_int16_d1[13]}} & {in_dat_data27, in_dat_data26});
    in_dat_data_int16_12 = ({16{cfg_is_int16_d1[12]}} & {in_dat_data25, in_dat_data24});
    in_dat_data_int16_11 = ({16{cfg_is_int16_d1[11]}} & {in_dat_data23, in_dat_data22});
    in_dat_data_int16_10 = ({16{cfg_is_int16_d1[10]}} & {in_dat_data21, in_dat_data20});
    in_dat_data_int16_9 = ({16{cfg_is_int16_d1[9]}} & {in_dat_data19, in_dat_data18});
    in_dat_data_int16_8 = ({16{cfg_is_int16_d1[8]}} & {in_dat_data17, in_dat_data16});
    in_dat_data_int16_7 = ({16{cfg_is_int16_d1[7]}} & {in_dat_data15, in_dat_data14});
    in_dat_data_int16_6 = ({16{cfg_is_int16_d1[6]}} & {in_dat_data13, in_dat_data12});
    in_dat_data_int16_5 = ({16{cfg_is_int16_d1[5]}} & {in_dat_data11, in_dat_data10});
    in_dat_data_int16_4 = ({16{cfg_is_int16_d1[4]}} & {in_dat_data9, in_dat_data8});
    in_dat_data_int16_3 = ({16{cfg_is_int16_d1[3]}} & {in_dat_data7, in_dat_data6});
    in_dat_data_int16_2 = ({16{cfg_is_int16_d1[2]}} & {in_dat_data5, in_dat_data4});
    in_dat_data_int16_1 = ({16{cfg_is_int16_d1[1]}} & {in_dat_data3, in_dat_data2});
    in_dat_data_int16_0 = ({16{cfg_is_int16_d1[0]}} & {in_dat_data1, in_dat_data0});
end



always @(
  in_dat_data_int16_63
  or in_dat_data_int16_62
  or in_dat_data_int16_61
  or in_dat_data_int16_60
  or in_dat_data_int16_59
  or in_dat_data_int16_58
  or in_dat_data_int16_57
  or in_dat_data_int16_56
  or in_dat_data_int16_55
  or in_dat_data_int16_54
  or in_dat_data_int16_53
  or in_dat_data_int16_52
  or in_dat_data_int16_51
  or in_dat_data_int16_50
  or in_dat_data_int16_49
  or in_dat_data_int16_48
  or in_dat_data_int16_47
  or in_dat_data_int16_46
  or in_dat_data_int16_45
  or in_dat_data_int16_44
  or in_dat_data_int16_43
  or in_dat_data_int16_42
  or in_dat_data_int16_41
  or in_dat_data_int16_40
  or in_dat_data_int16_39
  or in_dat_data_int16_38
  or in_dat_data_int16_37
  or in_dat_data_int16_36
  or in_dat_data_int16_35
  or in_dat_data_int16_34
  or in_dat_data_int16_33
  or in_dat_data_int16_32
  or in_dat_data_int16_31
  or in_dat_data_int16_30
  or in_dat_data_int16_29
  or in_dat_data_int16_28
  or in_dat_data_int16_27
  or in_dat_data_int16_26
  or in_dat_data_int16_25
  or in_dat_data_int16_24
  or in_dat_data_int16_23
  or in_dat_data_int16_22
  or in_dat_data_int16_21
  or in_dat_data_int16_20
  or in_dat_data_int16_19
  or in_dat_data_int16_18
  or in_dat_data_int16_17
  or in_dat_data_int16_16
  or in_dat_data_int16_15
  or in_dat_data_int16_14
  or in_dat_data_int16_13
  or in_dat_data_int16_12
  or in_dat_data_int16_11
  or in_dat_data_int16_10
  or in_dat_data_int16_9
  or in_dat_data_int16_8
  or in_dat_data_int16_7
  or in_dat_data_int16_6
  or in_dat_data_int16_5
  or in_dat_data_int16_4
  or in_dat_data_int16_3
  or in_dat_data_int16_2
  or in_dat_data_int16_1
  or in_dat_data_int16_0
  ) begin
    in_dat_data_int16 = {in_dat_data_int16_63, in_dat_data_int16_62, in_dat_data_int16_61, in_dat_data_int16_60, in_dat_data_int16_59, in_dat_data_int16_58, in_dat_data_int16_57, in_dat_data_int16_56, in_dat_data_int16_55, in_dat_data_int16_54, in_dat_data_int16_53, in_dat_data_int16_52, in_dat_data_int16_51, in_dat_data_int16_50, in_dat_data_int16_49, in_dat_data_int16_48, in_dat_data_int16_47, in_dat_data_int16_46, in_dat_data_int16_45, in_dat_data_int16_44, in_dat_data_int16_43, in_dat_data_int16_42, in_dat_data_int16_41, in_dat_data_int16_40, in_dat_data_int16_39, in_dat_data_int16_38, in_dat_data_int16_37, in_dat_data_int16_36, in_dat_data_int16_35, in_dat_data_int16_34, in_dat_data_int16_33, in_dat_data_int16_32, in_dat_data_int16_31, in_dat_data_int16_30, in_dat_data_int16_29, in_dat_data_int16_28, in_dat_data_int16_27, in_dat_data_int16_26, in_dat_data_int16_25, in_dat_data_int16_24, in_dat_data_int16_23, in_dat_data_int16_22, in_dat_data_int16_21, in_dat_data_int16_20, in_dat_data_int16_19, in_dat_data_int16_18, in_dat_data_int16_17, in_dat_data_int16_16, in_dat_data_int16_15, in_dat_data_int16_14, in_dat_data_int16_13, in_dat_data_int16_12, in_dat_data_int16_11, in_dat_data_int16_10, in_dat_data_int16_9, in_dat_data_int16_8, in_dat_data_int16_7, in_dat_data_int16_6, in_dat_data_int16_5, in_dat_data_int16_4, in_dat_data_int16_3, in_dat_data_int16_2, in_dat_data_int16_1, in_dat_data_int16_0};
end

//////////////// in_dat_data_int8 ////////////////
always @(
  cfg_is_int8_d1
  or in_dat_data127
  or in_dat_data63
  or in_dat_data126
  or in_dat_data62
  or in_dat_data125
  or in_dat_data61
  or in_dat_data124
  or in_dat_data60
  or in_dat_data123
  or in_dat_data59
  or in_dat_data122
  or in_dat_data58
  or in_dat_data121
  or in_dat_data57
  or in_dat_data120
  or in_dat_data56
  or in_dat_data119
  or in_dat_data55
  or in_dat_data118
  or in_dat_data54
  or in_dat_data117
  or in_dat_data53
  or in_dat_data116
  or in_dat_data52
  or in_dat_data115
  or in_dat_data51
  or in_dat_data114
  or in_dat_data50
  or in_dat_data113
  or in_dat_data49
  or in_dat_data112
  or in_dat_data48
  or in_dat_data111
  or in_dat_data47
  or in_dat_data110
  or in_dat_data46
  or in_dat_data109
  or in_dat_data45
  or in_dat_data108
  or in_dat_data44
  or in_dat_data107
  or in_dat_data43
  or in_dat_data106
  or in_dat_data42
  or in_dat_data105
  or in_dat_data41
  or in_dat_data104
  or in_dat_data40
  or in_dat_data103
  or in_dat_data39
  or in_dat_data102
  or in_dat_data38
  or in_dat_data101
  or in_dat_data37
  or in_dat_data100
  or in_dat_data36
  or in_dat_data99
  or in_dat_data35
  or in_dat_data98
  or in_dat_data34
  or in_dat_data97
  or in_dat_data33
  or in_dat_data96
  or in_dat_data32
  or in_dat_data95
  or in_dat_data31
  or in_dat_data94
  or in_dat_data30
  or in_dat_data93
  or in_dat_data29
  or in_dat_data92
  or in_dat_data28
  or in_dat_data91
  or in_dat_data27
  or in_dat_data90
  or in_dat_data26
  or in_dat_data89
  or in_dat_data25
  or in_dat_data88
  or in_dat_data24
  or in_dat_data87
  or in_dat_data23
  or in_dat_data86
  or in_dat_data22
  or in_dat_data85
  or in_dat_data21
  or in_dat_data84
  or in_dat_data20
  or in_dat_data83
  or in_dat_data19
  or in_dat_data82
  or in_dat_data18
  or in_dat_data81
  or in_dat_data17
  or in_dat_data80
  or in_dat_data16
  or in_dat_data79
  or in_dat_data15
  or in_dat_data78
  or in_dat_data14
  or in_dat_data77
  or in_dat_data13
  or in_dat_data76
  or in_dat_data12
  or in_dat_data75
  or in_dat_data11
  or in_dat_data74
  or in_dat_data10
  or in_dat_data73
  or in_dat_data9
  or in_dat_data72
  or in_dat_data8
  or in_dat_data71
  or in_dat_data7
  or in_dat_data70
  or in_dat_data6
  or in_dat_data69
  or in_dat_data5
  or in_dat_data68
  or in_dat_data4
  or in_dat_data67
  or in_dat_data3
  or in_dat_data66
  or in_dat_data2
  or in_dat_data65
  or in_dat_data1
  or in_dat_data64
  or in_dat_data0
  ) begin
    in_dat_data_int8_63 = ({16{cfg_is_int8_d1[63]}} & {in_dat_data127, in_dat_data63});
    in_dat_data_int8_62 = ({16{cfg_is_int8_d1[62]}} & {in_dat_data126, in_dat_data62});
    in_dat_data_int8_61 = ({16{cfg_is_int8_d1[61]}} & {in_dat_data125, in_dat_data61});
    in_dat_data_int8_60 = ({16{cfg_is_int8_d1[60]}} & {in_dat_data124, in_dat_data60});
    in_dat_data_int8_59 = ({16{cfg_is_int8_d1[59]}} & {in_dat_data123, in_dat_data59});
    in_dat_data_int8_58 = ({16{cfg_is_int8_d1[58]}} & {in_dat_data122, in_dat_data58});
    in_dat_data_int8_57 = ({16{cfg_is_int8_d1[57]}} & {in_dat_data121, in_dat_data57});
    in_dat_data_int8_56 = ({16{cfg_is_int8_d1[56]}} & {in_dat_data120, in_dat_data56});
    in_dat_data_int8_55 = ({16{cfg_is_int8_d1[55]}} & {in_dat_data119, in_dat_data55});
    in_dat_data_int8_54 = ({16{cfg_is_int8_d1[54]}} & {in_dat_data118, in_dat_data54});
    in_dat_data_int8_53 = ({16{cfg_is_int8_d1[53]}} & {in_dat_data117, in_dat_data53});
    in_dat_data_int8_52 = ({16{cfg_is_int8_d1[52]}} & {in_dat_data116, in_dat_data52});
    in_dat_data_int8_51 = ({16{cfg_is_int8_d1[51]}} & {in_dat_data115, in_dat_data51});
    in_dat_data_int8_50 = ({16{cfg_is_int8_d1[50]}} & {in_dat_data114, in_dat_data50});
    in_dat_data_int8_49 = ({16{cfg_is_int8_d1[49]}} & {in_dat_data113, in_dat_data49});
    in_dat_data_int8_48 = ({16{cfg_is_int8_d1[48]}} & {in_dat_data112, in_dat_data48});
    in_dat_data_int8_47 = ({16{cfg_is_int8_d1[47]}} & {in_dat_data111, in_dat_data47});
    in_dat_data_int8_46 = ({16{cfg_is_int8_d1[46]}} & {in_dat_data110, in_dat_data46});
    in_dat_data_int8_45 = ({16{cfg_is_int8_d1[45]}} & {in_dat_data109, in_dat_data45});
    in_dat_data_int8_44 = ({16{cfg_is_int8_d1[44]}} & {in_dat_data108, in_dat_data44});
    in_dat_data_int8_43 = ({16{cfg_is_int8_d1[43]}} & {in_dat_data107, in_dat_data43});
    in_dat_data_int8_42 = ({16{cfg_is_int8_d1[42]}} & {in_dat_data106, in_dat_data42});
    in_dat_data_int8_41 = ({16{cfg_is_int8_d1[41]}} & {in_dat_data105, in_dat_data41});
    in_dat_data_int8_40 = ({16{cfg_is_int8_d1[40]}} & {in_dat_data104, in_dat_data40});
    in_dat_data_int8_39 = ({16{cfg_is_int8_d1[39]}} & {in_dat_data103, in_dat_data39});
    in_dat_data_int8_38 = ({16{cfg_is_int8_d1[38]}} & {in_dat_data102, in_dat_data38});
    in_dat_data_int8_37 = ({16{cfg_is_int8_d1[37]}} & {in_dat_data101, in_dat_data37});
    in_dat_data_int8_36 = ({16{cfg_is_int8_d1[36]}} & {in_dat_data100, in_dat_data36});
    in_dat_data_int8_35 = ({16{cfg_is_int8_d1[35]}} & {in_dat_data99, in_dat_data35});
    in_dat_data_int8_34 = ({16{cfg_is_int8_d1[34]}} & {in_dat_data98, in_dat_data34});
    in_dat_data_int8_33 = ({16{cfg_is_int8_d1[33]}} & {in_dat_data97, in_dat_data33});
    in_dat_data_int8_32 = ({16{cfg_is_int8_d1[32]}} & {in_dat_data96, in_dat_data32});
    in_dat_data_int8_31 = ({16{cfg_is_int8_d1[31]}} & {in_dat_data95, in_dat_data31});
    in_dat_data_int8_30 = ({16{cfg_is_int8_d1[30]}} & {in_dat_data94, in_dat_data30});
    in_dat_data_int8_29 = ({16{cfg_is_int8_d1[29]}} & {in_dat_data93, in_dat_data29});
    in_dat_data_int8_28 = ({16{cfg_is_int8_d1[28]}} & {in_dat_data92, in_dat_data28});
    in_dat_data_int8_27 = ({16{cfg_is_int8_d1[27]}} & {in_dat_data91, in_dat_data27});
    in_dat_data_int8_26 = ({16{cfg_is_int8_d1[26]}} & {in_dat_data90, in_dat_data26});
    in_dat_data_int8_25 = ({16{cfg_is_int8_d1[25]}} & {in_dat_data89, in_dat_data25});
    in_dat_data_int8_24 = ({16{cfg_is_int8_d1[24]}} & {in_dat_data88, in_dat_data24});
    in_dat_data_int8_23 = ({16{cfg_is_int8_d1[23]}} & {in_dat_data87, in_dat_data23});
    in_dat_data_int8_22 = ({16{cfg_is_int8_d1[22]}} & {in_dat_data86, in_dat_data22});
    in_dat_data_int8_21 = ({16{cfg_is_int8_d1[21]}} & {in_dat_data85, in_dat_data21});
    in_dat_data_int8_20 = ({16{cfg_is_int8_d1[20]}} & {in_dat_data84, in_dat_data20});
    in_dat_data_int8_19 = ({16{cfg_is_int8_d1[19]}} & {in_dat_data83, in_dat_data19});
    in_dat_data_int8_18 = ({16{cfg_is_int8_d1[18]}} & {in_dat_data82, in_dat_data18});
    in_dat_data_int8_17 = ({16{cfg_is_int8_d1[17]}} & {in_dat_data81, in_dat_data17});
    in_dat_data_int8_16 = ({16{cfg_is_int8_d1[16]}} & {in_dat_data80, in_dat_data16});
    in_dat_data_int8_15 = ({16{cfg_is_int8_d1[15]}} & {in_dat_data79, in_dat_data15});
    in_dat_data_int8_14 = ({16{cfg_is_int8_d1[14]}} & {in_dat_data78, in_dat_data14});
    in_dat_data_int8_13 = ({16{cfg_is_int8_d1[13]}} & {in_dat_data77, in_dat_data13});
    in_dat_data_int8_12 = ({16{cfg_is_int8_d1[12]}} & {in_dat_data76, in_dat_data12});
    in_dat_data_int8_11 = ({16{cfg_is_int8_d1[11]}} & {in_dat_data75, in_dat_data11});
    in_dat_data_int8_10 = ({16{cfg_is_int8_d1[10]}} & {in_dat_data74, in_dat_data10});
    in_dat_data_int8_9 = ({16{cfg_is_int8_d1[9]}} & {in_dat_data73, in_dat_data9});
    in_dat_data_int8_8 = ({16{cfg_is_int8_d1[8]}} & {in_dat_data72, in_dat_data8});
    in_dat_data_int8_7 = ({16{cfg_is_int8_d1[7]}} & {in_dat_data71, in_dat_data7});
    in_dat_data_int8_6 = ({16{cfg_is_int8_d1[6]}} & {in_dat_data70, in_dat_data6});
    in_dat_data_int8_5 = ({16{cfg_is_int8_d1[5]}} & {in_dat_data69, in_dat_data5});
    in_dat_data_int8_4 = ({16{cfg_is_int8_d1[4]}} & {in_dat_data68, in_dat_data4});
    in_dat_data_int8_3 = ({16{cfg_is_int8_d1[3]}} & {in_dat_data67, in_dat_data3});
    in_dat_data_int8_2 = ({16{cfg_is_int8_d1[2]}} & {in_dat_data66, in_dat_data2});
    in_dat_data_int8_1 = ({16{cfg_is_int8_d1[1]}} & {in_dat_data65, in_dat_data1});
    in_dat_data_int8_0 = ({16{cfg_is_int8_d1[0]}} & {in_dat_data64, in_dat_data0});
end


always @(
  in_dat_mask
  ) begin
    in_dat_mask_int8 = {in_dat_mask[127], in_dat_mask[63], in_dat_mask[126], in_dat_mask[62], in_dat_mask[125], in_dat_mask[61], in_dat_mask[124], in_dat_mask[60], in_dat_mask[123], in_dat_mask[59], in_dat_mask[122], in_dat_mask[58], in_dat_mask[121], in_dat_mask[57], in_dat_mask[120], in_dat_mask[56],
                        in_dat_mask[119], in_dat_mask[55], in_dat_mask[118], in_dat_mask[54], in_dat_mask[117], in_dat_mask[53], in_dat_mask[116], in_dat_mask[52], in_dat_mask[115], in_dat_mask[51], in_dat_mask[114], in_dat_mask[50], in_dat_mask[113], in_dat_mask[49], in_dat_mask[112], in_dat_mask[48],
                        in_dat_mask[111], in_dat_mask[47], in_dat_mask[110], in_dat_mask[46], in_dat_mask[109], in_dat_mask[45], in_dat_mask[108], in_dat_mask[44], in_dat_mask[107], in_dat_mask[43], in_dat_mask[106], in_dat_mask[42], in_dat_mask[105], in_dat_mask[41], in_dat_mask[104], in_dat_mask[40],
                        in_dat_mask[103], in_dat_mask[39], in_dat_mask[102], in_dat_mask[38], in_dat_mask[101], in_dat_mask[37], in_dat_mask[100], in_dat_mask[36], in_dat_mask[99], in_dat_mask[35], in_dat_mask[98], in_dat_mask[34], in_dat_mask[97], in_dat_mask[33], in_dat_mask[96], in_dat_mask[32],
                        in_dat_mask[95], in_dat_mask[31], in_dat_mask[94], in_dat_mask[30], in_dat_mask[93], in_dat_mask[29], in_dat_mask[92], in_dat_mask[28], in_dat_mask[91], in_dat_mask[27], in_dat_mask[90], in_dat_mask[26], in_dat_mask[89], in_dat_mask[25], in_dat_mask[88], in_dat_mask[24],
                        in_dat_mask[87], in_dat_mask[23], in_dat_mask[86], in_dat_mask[22], in_dat_mask[85], in_dat_mask[21], in_dat_mask[84], in_dat_mask[20], in_dat_mask[83], in_dat_mask[19], in_dat_mask[82], in_dat_mask[18], in_dat_mask[81], in_dat_mask[17], in_dat_mask[80], in_dat_mask[16],
                        in_dat_mask[79], in_dat_mask[15], in_dat_mask[78], in_dat_mask[14], in_dat_mask[77], in_dat_mask[13], in_dat_mask[76], in_dat_mask[12], in_dat_mask[75], in_dat_mask[11], in_dat_mask[74], in_dat_mask[10], in_dat_mask[73], in_dat_mask[9], in_dat_mask[72], in_dat_mask[8],
                        in_dat_mask[71], in_dat_mask[7], in_dat_mask[70], in_dat_mask[6], in_dat_mask[69], in_dat_mask[5], in_dat_mask[68], in_dat_mask[4], in_dat_mask[67], in_dat_mask[3], in_dat_mask[66], in_dat_mask[2], in_dat_mask[65], in_dat_mask[1], in_dat_mask[64], in_dat_mask[0]};
end



always @(
  in_dat_data_int8_63
  or in_dat_data_int8_62
  or in_dat_data_int8_61
  or in_dat_data_int8_60
  or in_dat_data_int8_59
  or in_dat_data_int8_58
  or in_dat_data_int8_57
  or in_dat_data_int8_56
  or in_dat_data_int8_55
  or in_dat_data_int8_54
  or in_dat_data_int8_53
  or in_dat_data_int8_52
  or in_dat_data_int8_51
  or in_dat_data_int8_50
  or in_dat_data_int8_49
  or in_dat_data_int8_48
  or in_dat_data_int8_47
  or in_dat_data_int8_46
  or in_dat_data_int8_45
  or in_dat_data_int8_44
  or in_dat_data_int8_43
  or in_dat_data_int8_42
  or in_dat_data_int8_41
  or in_dat_data_int8_40
  or in_dat_data_int8_39
  or in_dat_data_int8_38
  or in_dat_data_int8_37
  or in_dat_data_int8_36
  or in_dat_data_int8_35
  or in_dat_data_int8_34
  or in_dat_data_int8_33
  or in_dat_data_int8_32
  or in_dat_data_int8_31
  or in_dat_data_int8_30
  or in_dat_data_int8_29
  or in_dat_data_int8_28
  or in_dat_data_int8_27
  or in_dat_data_int8_26
  or in_dat_data_int8_25
  or in_dat_data_int8_24
  or in_dat_data_int8_23
  or in_dat_data_int8_22
  or in_dat_data_int8_21
  or in_dat_data_int8_20
  or in_dat_data_int8_19
  or in_dat_data_int8_18
  or in_dat_data_int8_17
  or in_dat_data_int8_16
  or in_dat_data_int8_15
  or in_dat_data_int8_14
  or in_dat_data_int8_13
  or in_dat_data_int8_12
  or in_dat_data_int8_11
  or in_dat_data_int8_10
  or in_dat_data_int8_9
  or in_dat_data_int8_8
  or in_dat_data_int8_7
  or in_dat_data_int8_6
  or in_dat_data_int8_5
  or in_dat_data_int8_4
  or in_dat_data_int8_3
  or in_dat_data_int8_2
  or in_dat_data_int8_1
  or in_dat_data_int8_0
  ) begin
    in_dat_data_int8 = {in_dat_data_int8_63, in_dat_data_int8_62, in_dat_data_int8_61, in_dat_data_int8_60, in_dat_data_int8_59, in_dat_data_int8_58, in_dat_data_int8_57, in_dat_data_int8_56, in_dat_data_int8_55, in_dat_data_int8_54, in_dat_data_int8_53, in_dat_data_int8_52, in_dat_data_int8_51, in_dat_data_int8_50, in_dat_data_int8_49, in_dat_data_int8_48, in_dat_data_int8_47, in_dat_data_int8_46, in_dat_data_int8_45, in_dat_data_int8_44, in_dat_data_int8_43, in_dat_data_int8_42, in_dat_data_int8_41, in_dat_data_int8_40, in_dat_data_int8_39, in_dat_data_int8_38, in_dat_data_int8_37, in_dat_data_int8_36, in_dat_data_int8_35, in_dat_data_int8_34, in_dat_data_int8_33, in_dat_data_int8_32, in_dat_data_int8_31, in_dat_data_int8_30, in_dat_data_int8_29, in_dat_data_int8_28, in_dat_data_int8_27, in_dat_data_int8_26, in_dat_data_int8_25, in_dat_data_int8_24, in_dat_data_int8_23, in_dat_data_int8_22, in_dat_data_int8_21, in_dat_data_int8_20, in_dat_data_int8_19, in_dat_data_int8_18, in_dat_data_int8_17, in_dat_data_int8_16, in_dat_data_int8_15, in_dat_data_int8_14, in_dat_data_int8_13, in_dat_data_int8_12, in_dat_data_int8_11, in_dat_data_int8_10, in_dat_data_int8_9, in_dat_data_int8_8, in_dat_data_int8_7, in_dat_data_int8_6, in_dat_data_int8_5, in_dat_data_int8_4, in_dat_data_int8_3, in_dat_data_int8_2, in_dat_data_int8_1, in_dat_data_int8_0};
end

//////////////// in_dat_data_fp16 ////////////////

always @(
  cfg_is_fp16_d1
  or in_dat_data_pack
  or in_dat_mask
  ) begin
    in_dat_nan[63] = cfg_is_fp16_d1[63] & (&in_dat_data_pack[1022:1018]) & (|in_dat_data_pack[1017:1008]) & in_dat_mask[126];
    in_dat_nan[62] = cfg_is_fp16_d1[62] & (&in_dat_data_pack[1006:1002]) & (|in_dat_data_pack[1001:992]) & in_dat_mask[124];
    in_dat_nan[61] = cfg_is_fp16_d1[61] & (&in_dat_data_pack[990:986]) & (|in_dat_data_pack[985:976]) & in_dat_mask[122];
    in_dat_nan[60] = cfg_is_fp16_d1[60] & (&in_dat_data_pack[974:970]) & (|in_dat_data_pack[969:960]) & in_dat_mask[120];
    in_dat_nan[59] = cfg_is_fp16_d1[59] & (&in_dat_data_pack[958:954]) & (|in_dat_data_pack[953:944]) & in_dat_mask[118];
    in_dat_nan[58] = cfg_is_fp16_d1[58] & (&in_dat_data_pack[942:938]) & (|in_dat_data_pack[937:928]) & in_dat_mask[116];
    in_dat_nan[57] = cfg_is_fp16_d1[57] & (&in_dat_data_pack[926:922]) & (|in_dat_data_pack[921:912]) & in_dat_mask[114];
    in_dat_nan[56] = cfg_is_fp16_d1[56] & (&in_dat_data_pack[910:906]) & (|in_dat_data_pack[905:896]) & in_dat_mask[112];
    in_dat_nan[55] = cfg_is_fp16_d1[55] & (&in_dat_data_pack[894:890]) & (|in_dat_data_pack[889:880]) & in_dat_mask[110];
    in_dat_nan[54] = cfg_is_fp16_d1[54] & (&in_dat_data_pack[878:874]) & (|in_dat_data_pack[873:864]) & in_dat_mask[108];
    in_dat_nan[53] = cfg_is_fp16_d1[53] & (&in_dat_data_pack[862:858]) & (|in_dat_data_pack[857:848]) & in_dat_mask[106];
    in_dat_nan[52] = cfg_is_fp16_d1[52] & (&in_dat_data_pack[846:842]) & (|in_dat_data_pack[841:832]) & in_dat_mask[104];
    in_dat_nan[51] = cfg_is_fp16_d1[51] & (&in_dat_data_pack[830:826]) & (|in_dat_data_pack[825:816]) & in_dat_mask[102];
    in_dat_nan[50] = cfg_is_fp16_d1[50] & (&in_dat_data_pack[814:810]) & (|in_dat_data_pack[809:800]) & in_dat_mask[100];
    in_dat_nan[49] = cfg_is_fp16_d1[49] & (&in_dat_data_pack[798:794]) & (|in_dat_data_pack[793:784]) & in_dat_mask[98];
    in_dat_nan[48] = cfg_is_fp16_d1[48] & (&in_dat_data_pack[782:778]) & (|in_dat_data_pack[777:768]) & in_dat_mask[96];
    in_dat_nan[47] = cfg_is_fp16_d1[47] & (&in_dat_data_pack[766:762]) & (|in_dat_data_pack[761:752]) & in_dat_mask[94];
    in_dat_nan[46] = cfg_is_fp16_d1[46] & (&in_dat_data_pack[750:746]) & (|in_dat_data_pack[745:736]) & in_dat_mask[92];
    in_dat_nan[45] = cfg_is_fp16_d1[45] & (&in_dat_data_pack[734:730]) & (|in_dat_data_pack[729:720]) & in_dat_mask[90];
    in_dat_nan[44] = cfg_is_fp16_d1[44] & (&in_dat_data_pack[718:714]) & (|in_dat_data_pack[713:704]) & in_dat_mask[88];
    in_dat_nan[43] = cfg_is_fp16_d1[43] & (&in_dat_data_pack[702:698]) & (|in_dat_data_pack[697:688]) & in_dat_mask[86];
    in_dat_nan[42] = cfg_is_fp16_d1[42] & (&in_dat_data_pack[686:682]) & (|in_dat_data_pack[681:672]) & in_dat_mask[84];
    in_dat_nan[41] = cfg_is_fp16_d1[41] & (&in_dat_data_pack[670:666]) & (|in_dat_data_pack[665:656]) & in_dat_mask[82];
    in_dat_nan[40] = cfg_is_fp16_d1[40] & (&in_dat_data_pack[654:650]) & (|in_dat_data_pack[649:640]) & in_dat_mask[80];
    in_dat_nan[39] = cfg_is_fp16_d1[39] & (&in_dat_data_pack[638:634]) & (|in_dat_data_pack[633:624]) & in_dat_mask[78];
    in_dat_nan[38] = cfg_is_fp16_d1[38] & (&in_dat_data_pack[622:618]) & (|in_dat_data_pack[617:608]) & in_dat_mask[76];
    in_dat_nan[37] = cfg_is_fp16_d1[37] & (&in_dat_data_pack[606:602]) & (|in_dat_data_pack[601:592]) & in_dat_mask[74];
    in_dat_nan[36] = cfg_is_fp16_d1[36] & (&in_dat_data_pack[590:586]) & (|in_dat_data_pack[585:576]) & in_dat_mask[72];
    in_dat_nan[35] = cfg_is_fp16_d1[35] & (&in_dat_data_pack[574:570]) & (|in_dat_data_pack[569:560]) & in_dat_mask[70];
    in_dat_nan[34] = cfg_is_fp16_d1[34] & (&in_dat_data_pack[558:554]) & (|in_dat_data_pack[553:544]) & in_dat_mask[68];
    in_dat_nan[33] = cfg_is_fp16_d1[33] & (&in_dat_data_pack[542:538]) & (|in_dat_data_pack[537:528]) & in_dat_mask[66];
    in_dat_nan[32] = cfg_is_fp16_d1[32] & (&in_dat_data_pack[526:522]) & (|in_dat_data_pack[521:512]) & in_dat_mask[64];
    in_dat_nan[31] = cfg_is_fp16_d1[31] & (&in_dat_data_pack[510:506]) & (|in_dat_data_pack[505:496]) & in_dat_mask[62];
    in_dat_nan[30] = cfg_is_fp16_d1[30] & (&in_dat_data_pack[494:490]) & (|in_dat_data_pack[489:480]) & in_dat_mask[60];
    in_dat_nan[29] = cfg_is_fp16_d1[29] & (&in_dat_data_pack[478:474]) & (|in_dat_data_pack[473:464]) & in_dat_mask[58];
    in_dat_nan[28] = cfg_is_fp16_d1[28] & (&in_dat_data_pack[462:458]) & (|in_dat_data_pack[457:448]) & in_dat_mask[56];
    in_dat_nan[27] = cfg_is_fp16_d1[27] & (&in_dat_data_pack[446:442]) & (|in_dat_data_pack[441:432]) & in_dat_mask[54];
    in_dat_nan[26] = cfg_is_fp16_d1[26] & (&in_dat_data_pack[430:426]) & (|in_dat_data_pack[425:416]) & in_dat_mask[52];
    in_dat_nan[25] = cfg_is_fp16_d1[25] & (&in_dat_data_pack[414:410]) & (|in_dat_data_pack[409:400]) & in_dat_mask[50];
    in_dat_nan[24] = cfg_is_fp16_d1[24] & (&in_dat_data_pack[398:394]) & (|in_dat_data_pack[393:384]) & in_dat_mask[48];
    in_dat_nan[23] = cfg_is_fp16_d1[23] & (&in_dat_data_pack[382:378]) & (|in_dat_data_pack[377:368]) & in_dat_mask[46];
    in_dat_nan[22] = cfg_is_fp16_d1[22] & (&in_dat_data_pack[366:362]) & (|in_dat_data_pack[361:352]) & in_dat_mask[44];
    in_dat_nan[21] = cfg_is_fp16_d1[21] & (&in_dat_data_pack[350:346]) & (|in_dat_data_pack[345:336]) & in_dat_mask[42];
    in_dat_nan[20] = cfg_is_fp16_d1[20] & (&in_dat_data_pack[334:330]) & (|in_dat_data_pack[329:320]) & in_dat_mask[40];
    in_dat_nan[19] = cfg_is_fp16_d1[19] & (&in_dat_data_pack[318:314]) & (|in_dat_data_pack[313:304]) & in_dat_mask[38];
    in_dat_nan[18] = cfg_is_fp16_d1[18] & (&in_dat_data_pack[302:298]) & (|in_dat_data_pack[297:288]) & in_dat_mask[36];
    in_dat_nan[17] = cfg_is_fp16_d1[17] & (&in_dat_data_pack[286:282]) & (|in_dat_data_pack[281:272]) & in_dat_mask[34];
    in_dat_nan[16] = cfg_is_fp16_d1[16] & (&in_dat_data_pack[270:266]) & (|in_dat_data_pack[265:256]) & in_dat_mask[32];
    in_dat_nan[15] = cfg_is_fp16_d1[15] & (&in_dat_data_pack[254:250]) & (|in_dat_data_pack[249:240]) & in_dat_mask[30];
    in_dat_nan[14] = cfg_is_fp16_d1[14] & (&in_dat_data_pack[238:234]) & (|in_dat_data_pack[233:224]) & in_dat_mask[28];
    in_dat_nan[13] = cfg_is_fp16_d1[13] & (&in_dat_data_pack[222:218]) & (|in_dat_data_pack[217:208]) & in_dat_mask[26];
    in_dat_nan[12] = cfg_is_fp16_d1[12] & (&in_dat_data_pack[206:202]) & (|in_dat_data_pack[201:192]) & in_dat_mask[24];
    in_dat_nan[11] = cfg_is_fp16_d1[11] & (&in_dat_data_pack[190:186]) & (|in_dat_data_pack[185:176]) & in_dat_mask[22];
    in_dat_nan[10] = cfg_is_fp16_d1[10] & (&in_dat_data_pack[174:170]) & (|in_dat_data_pack[169:160]) & in_dat_mask[20];
    in_dat_nan[9] = cfg_is_fp16_d1[9] & (&in_dat_data_pack[158:154]) & (|in_dat_data_pack[153:144]) & in_dat_mask[18];
    in_dat_nan[8] = cfg_is_fp16_d1[8] & (&in_dat_data_pack[142:138]) & (|in_dat_data_pack[137:128]) & in_dat_mask[16];
    in_dat_nan[7] = cfg_is_fp16_d1[7] & (&in_dat_data_pack[126:122]) & (|in_dat_data_pack[121:112]) & in_dat_mask[14];
    in_dat_nan[6] = cfg_is_fp16_d1[6] & (&in_dat_data_pack[110:106]) & (|in_dat_data_pack[105:96]) & in_dat_mask[12];
    in_dat_nan[5] = cfg_is_fp16_d1[5] & (&in_dat_data_pack[94:90]) & (|in_dat_data_pack[89:80]) & in_dat_mask[10];
    in_dat_nan[4] = cfg_is_fp16_d1[4] & (&in_dat_data_pack[78:74]) & (|in_dat_data_pack[73:64]) & in_dat_mask[8];
    in_dat_nan[3] = cfg_is_fp16_d1[3] & (&in_dat_data_pack[62:58]) & (|in_dat_data_pack[57:48]) & in_dat_mask[6];
    in_dat_nan[2] = cfg_is_fp16_d1[2] & (&in_dat_data_pack[46:42]) & (|in_dat_data_pack[41:32]) & in_dat_mask[4];
    in_dat_nan[1] = cfg_is_fp16_d1[1] & (&in_dat_data_pack[30:26]) & (|in_dat_data_pack[25:16]) & in_dat_mask[2];
    in_dat_nan[0] = cfg_is_fp16_d1[0] & (&in_dat_data_pack[14:10]) & (|in_dat_data_pack[9:0]) & in_dat_mask[0];
end


always @(
  cfg_is_fp16_d1
  or in_dat_mask
  or in_dat_data_pack
  ) begin
    in_dat_exp[191:189] = {3{cfg_is_fp16_d1[63] & in_dat_mask[127]}} & (in_dat_data_pack[1022:1020]);
    in_dat_exp[188:186] = {3{cfg_is_fp16_d1[62] & in_dat_mask[125]}} & (in_dat_data_pack[1006:1004]);
    in_dat_exp[185:183] = {3{cfg_is_fp16_d1[61] & in_dat_mask[123]}} & (in_dat_data_pack[990:988]);
    in_dat_exp[182:180] = {3{cfg_is_fp16_d1[60] & in_dat_mask[121]}} & (in_dat_data_pack[974:972]);
    in_dat_exp[179:177] = {3{cfg_is_fp16_d1[59] & in_dat_mask[119]}} & (in_dat_data_pack[958:956]);
    in_dat_exp[176:174] = {3{cfg_is_fp16_d1[58] & in_dat_mask[117]}} & (in_dat_data_pack[942:940]);
    in_dat_exp[173:171] = {3{cfg_is_fp16_d1[57] & in_dat_mask[115]}} & (in_dat_data_pack[926:924]);
    in_dat_exp[170:168] = {3{cfg_is_fp16_d1[56] & in_dat_mask[113]}} & (in_dat_data_pack[910:908]);
    in_dat_exp[167:165] = {3{cfg_is_fp16_d1[55] & in_dat_mask[111]}} & (in_dat_data_pack[894:892]);
    in_dat_exp[164:162] = {3{cfg_is_fp16_d1[54] & in_dat_mask[109]}} & (in_dat_data_pack[878:876]);
    in_dat_exp[161:159] = {3{cfg_is_fp16_d1[53] & in_dat_mask[107]}} & (in_dat_data_pack[862:860]);
    in_dat_exp[158:156] = {3{cfg_is_fp16_d1[52] & in_dat_mask[105]}} & (in_dat_data_pack[846:844]);
    in_dat_exp[155:153] = {3{cfg_is_fp16_d1[51] & in_dat_mask[103]}} & (in_dat_data_pack[830:828]);
    in_dat_exp[152:150] = {3{cfg_is_fp16_d1[50] & in_dat_mask[101]}} & (in_dat_data_pack[814:812]);
    in_dat_exp[149:147] = {3{cfg_is_fp16_d1[49] & in_dat_mask[99]}} & (in_dat_data_pack[798:796]);
    in_dat_exp[146:144] = {3{cfg_is_fp16_d1[48] & in_dat_mask[97]}} & (in_dat_data_pack[782:780]);
    in_dat_exp[143:141] = {3{cfg_is_fp16_d1[47] & in_dat_mask[95]}} & (in_dat_data_pack[766:764]);
    in_dat_exp[140:138] = {3{cfg_is_fp16_d1[46] & in_dat_mask[93]}} & (in_dat_data_pack[750:748]);
    in_dat_exp[137:135] = {3{cfg_is_fp16_d1[45] & in_dat_mask[91]}} & (in_dat_data_pack[734:732]);
    in_dat_exp[134:132] = {3{cfg_is_fp16_d1[44] & in_dat_mask[89]}} & (in_dat_data_pack[718:716]);
    in_dat_exp[131:129] = {3{cfg_is_fp16_d1[43] & in_dat_mask[87]}} & (in_dat_data_pack[702:700]);
    in_dat_exp[128:126] = {3{cfg_is_fp16_d1[42] & in_dat_mask[85]}} & (in_dat_data_pack[686:684]);
    in_dat_exp[125:123] = {3{cfg_is_fp16_d1[41] & in_dat_mask[83]}} & (in_dat_data_pack[670:668]);
    in_dat_exp[122:120] = {3{cfg_is_fp16_d1[40] & in_dat_mask[81]}} & (in_dat_data_pack[654:652]);
    in_dat_exp[119:117] = {3{cfg_is_fp16_d1[39] & in_dat_mask[79]}} & (in_dat_data_pack[638:636]);
    in_dat_exp[116:114] = {3{cfg_is_fp16_d1[38] & in_dat_mask[77]}} & (in_dat_data_pack[622:620]);
    in_dat_exp[113:111] = {3{cfg_is_fp16_d1[37] & in_dat_mask[75]}} & (in_dat_data_pack[606:604]);
    in_dat_exp[110:108] = {3{cfg_is_fp16_d1[36] & in_dat_mask[73]}} & (in_dat_data_pack[590:588]);
    in_dat_exp[107:105] = {3{cfg_is_fp16_d1[35] & in_dat_mask[71]}} & (in_dat_data_pack[574:572]);
    in_dat_exp[104:102] = {3{cfg_is_fp16_d1[34] & in_dat_mask[69]}} & (in_dat_data_pack[558:556]);
    in_dat_exp[101:99] = {3{cfg_is_fp16_d1[33] & in_dat_mask[67]}} & (in_dat_data_pack[542:540]);
    in_dat_exp[98:96] = {3{cfg_is_fp16_d1[32] & in_dat_mask[65]}} & (in_dat_data_pack[526:524]);
    in_dat_exp[95:93] = {3{cfg_is_fp16_d1[31] & in_dat_mask[63]}} & (in_dat_data_pack[510:508]);
    in_dat_exp[92:90] = {3{cfg_is_fp16_d1[30] & in_dat_mask[61]}} & (in_dat_data_pack[494:492]);
    in_dat_exp[89:87] = {3{cfg_is_fp16_d1[29] & in_dat_mask[59]}} & (in_dat_data_pack[478:476]);
    in_dat_exp[86:84] = {3{cfg_is_fp16_d1[28] & in_dat_mask[57]}} & (in_dat_data_pack[462:460]);
    in_dat_exp[83:81] = {3{cfg_is_fp16_d1[27] & in_dat_mask[55]}} & (in_dat_data_pack[446:444]);
    in_dat_exp[80:78] = {3{cfg_is_fp16_d1[26] & in_dat_mask[53]}} & (in_dat_data_pack[430:428]);
    in_dat_exp[77:75] = {3{cfg_is_fp16_d1[25] & in_dat_mask[51]}} & (in_dat_data_pack[414:412]);
    in_dat_exp[74:72] = {3{cfg_is_fp16_d1[24] & in_dat_mask[49]}} & (in_dat_data_pack[398:396]);
    in_dat_exp[71:69] = {3{cfg_is_fp16_d1[23] & in_dat_mask[47]}} & (in_dat_data_pack[382:380]);
    in_dat_exp[68:66] = {3{cfg_is_fp16_d1[22] & in_dat_mask[45]}} & (in_dat_data_pack[366:364]);
    in_dat_exp[65:63] = {3{cfg_is_fp16_d1[21] & in_dat_mask[43]}} & (in_dat_data_pack[350:348]);
    in_dat_exp[62:60] = {3{cfg_is_fp16_d1[20] & in_dat_mask[41]}} & (in_dat_data_pack[334:332]);
    in_dat_exp[59:57] = {3{cfg_is_fp16_d1[19] & in_dat_mask[39]}} & (in_dat_data_pack[318:316]);
    in_dat_exp[56:54] = {3{cfg_is_fp16_d1[18] & in_dat_mask[37]}} & (in_dat_data_pack[302:300]);
    in_dat_exp[53:51] = {3{cfg_is_fp16_d1[17] & in_dat_mask[35]}} & (in_dat_data_pack[286:284]);
    in_dat_exp[50:48] = {3{cfg_is_fp16_d1[16] & in_dat_mask[33]}} & (in_dat_data_pack[270:268]);
    in_dat_exp[47:45] = {3{cfg_is_fp16_d1[15] & in_dat_mask[31]}} & (in_dat_data_pack[254:252]);
    in_dat_exp[44:42] = {3{cfg_is_fp16_d1[14] & in_dat_mask[29]}} & (in_dat_data_pack[238:236]);
    in_dat_exp[41:39] = {3{cfg_is_fp16_d1[13] & in_dat_mask[27]}} & (in_dat_data_pack[222:220]);
    in_dat_exp[38:36] = {3{cfg_is_fp16_d1[12] & in_dat_mask[25]}} & (in_dat_data_pack[206:204]);
    in_dat_exp[35:33] = {3{cfg_is_fp16_d1[11] & in_dat_mask[23]}} & (in_dat_data_pack[190:188]);
    in_dat_exp[32:30] = {3{cfg_is_fp16_d1[10] & in_dat_mask[21]}} & (in_dat_data_pack[174:172]);
    in_dat_exp[29:27] = {3{cfg_is_fp16_d1[9] & in_dat_mask[19]}} & (in_dat_data_pack[158:156]);
    in_dat_exp[26:24] = {3{cfg_is_fp16_d1[8] & in_dat_mask[17]}} & (in_dat_data_pack[142:140]);
    in_dat_exp[23:21] = {3{cfg_is_fp16_d1[7] & in_dat_mask[15]}} & (in_dat_data_pack[126:124]);
    in_dat_exp[20:18] = {3{cfg_is_fp16_d1[6] & in_dat_mask[13]}} & (in_dat_data_pack[110:108]);
    in_dat_exp[17:15] = {3{cfg_is_fp16_d1[5] & in_dat_mask[11]}} & (in_dat_data_pack[94:92]);
    in_dat_exp[14:12] = {3{cfg_is_fp16_d1[4] & in_dat_mask[9]}} & (in_dat_data_pack[78:76]);
    in_dat_exp[11:9] = {3{cfg_is_fp16_d1[3] & in_dat_mask[7]}} & (in_dat_data_pack[62:60]);
    in_dat_exp[8:6] = {3{cfg_is_fp16_d1[2] & in_dat_mask[5]}} & (in_dat_data_pack[46:44]);
    in_dat_exp[5:3] = {3{cfg_is_fp16_d1[1] & in_dat_mask[3]}} & (in_dat_data_pack[30:28]);
    in_dat_exp[2:0] = {3{cfg_is_fp16_d1[0] & in_dat_mask[1]}} & (in_dat_data_pack[14:12]);
end


always @(
  cfg_is_fp16_d1
  or in_dat_data_pack
  ) begin
    in_dat_norm[63] = cfg_is_fp16_d1[63] & (|in_dat_data_pack[1022:1018]);
    in_dat_norm[62] = cfg_is_fp16_d1[62] & (|in_dat_data_pack[1006:1002]);
    in_dat_norm[61] = cfg_is_fp16_d1[61] & (|in_dat_data_pack[990:986]);
    in_dat_norm[60] = cfg_is_fp16_d1[60] & (|in_dat_data_pack[974:970]);
    in_dat_norm[59] = cfg_is_fp16_d1[59] & (|in_dat_data_pack[958:954]);
    in_dat_norm[58] = cfg_is_fp16_d1[58] & (|in_dat_data_pack[942:938]);
    in_dat_norm[57] = cfg_is_fp16_d1[57] & (|in_dat_data_pack[926:922]);
    in_dat_norm[56] = cfg_is_fp16_d1[56] & (|in_dat_data_pack[910:906]);
    in_dat_norm[55] = cfg_is_fp16_d1[55] & (|in_dat_data_pack[894:890]);
    in_dat_norm[54] = cfg_is_fp16_d1[54] & (|in_dat_data_pack[878:874]);
    in_dat_norm[53] = cfg_is_fp16_d1[53] & (|in_dat_data_pack[862:858]);
    in_dat_norm[52] = cfg_is_fp16_d1[52] & (|in_dat_data_pack[846:842]);
    in_dat_norm[51] = cfg_is_fp16_d1[51] & (|in_dat_data_pack[830:826]);
    in_dat_norm[50] = cfg_is_fp16_d1[50] & (|in_dat_data_pack[814:810]);
    in_dat_norm[49] = cfg_is_fp16_d1[49] & (|in_dat_data_pack[798:794]);
    in_dat_norm[48] = cfg_is_fp16_d1[48] & (|in_dat_data_pack[782:778]);
    in_dat_norm[47] = cfg_is_fp16_d1[47] & (|in_dat_data_pack[766:762]);
    in_dat_norm[46] = cfg_is_fp16_d1[46] & (|in_dat_data_pack[750:746]);
    in_dat_norm[45] = cfg_is_fp16_d1[45] & (|in_dat_data_pack[734:730]);
    in_dat_norm[44] = cfg_is_fp16_d1[44] & (|in_dat_data_pack[718:714]);
    in_dat_norm[43] = cfg_is_fp16_d1[43] & (|in_dat_data_pack[702:698]);
    in_dat_norm[42] = cfg_is_fp16_d1[42] & (|in_dat_data_pack[686:682]);
    in_dat_norm[41] = cfg_is_fp16_d1[41] & (|in_dat_data_pack[670:666]);
    in_dat_norm[40] = cfg_is_fp16_d1[40] & (|in_dat_data_pack[654:650]);
    in_dat_norm[39] = cfg_is_fp16_d1[39] & (|in_dat_data_pack[638:634]);
    in_dat_norm[38] = cfg_is_fp16_d1[38] & (|in_dat_data_pack[622:618]);
    in_dat_norm[37] = cfg_is_fp16_d1[37] & (|in_dat_data_pack[606:602]);
    in_dat_norm[36] = cfg_is_fp16_d1[36] & (|in_dat_data_pack[590:586]);
    in_dat_norm[35] = cfg_is_fp16_d1[35] & (|in_dat_data_pack[574:570]);
    in_dat_norm[34] = cfg_is_fp16_d1[34] & (|in_dat_data_pack[558:554]);
    in_dat_norm[33] = cfg_is_fp16_d1[33] & (|in_dat_data_pack[542:538]);
    in_dat_norm[32] = cfg_is_fp16_d1[32] & (|in_dat_data_pack[526:522]);
    in_dat_norm[31] = cfg_is_fp16_d1[31] & (|in_dat_data_pack[510:506]);
    in_dat_norm[30] = cfg_is_fp16_d1[30] & (|in_dat_data_pack[494:490]);
    in_dat_norm[29] = cfg_is_fp16_d1[29] & (|in_dat_data_pack[478:474]);
    in_dat_norm[28] = cfg_is_fp16_d1[28] & (|in_dat_data_pack[462:458]);
    in_dat_norm[27] = cfg_is_fp16_d1[27] & (|in_dat_data_pack[446:442]);
    in_dat_norm[26] = cfg_is_fp16_d1[26] & (|in_dat_data_pack[430:426]);
    in_dat_norm[25] = cfg_is_fp16_d1[25] & (|in_dat_data_pack[414:410]);
    in_dat_norm[24] = cfg_is_fp16_d1[24] & (|in_dat_data_pack[398:394]);
    in_dat_norm[23] = cfg_is_fp16_d1[23] & (|in_dat_data_pack[382:378]);
    in_dat_norm[22] = cfg_is_fp16_d1[22] & (|in_dat_data_pack[366:362]);
    in_dat_norm[21] = cfg_is_fp16_d1[21] & (|in_dat_data_pack[350:346]);
    in_dat_norm[20] = cfg_is_fp16_d1[20] & (|in_dat_data_pack[334:330]);
    in_dat_norm[19] = cfg_is_fp16_d1[19] & (|in_dat_data_pack[318:314]);
    in_dat_norm[18] = cfg_is_fp16_d1[18] & (|in_dat_data_pack[302:298]);
    in_dat_norm[17] = cfg_is_fp16_d1[17] & (|in_dat_data_pack[286:282]);
    in_dat_norm[16] = cfg_is_fp16_d1[16] & (|in_dat_data_pack[270:266]);
    in_dat_norm[15] = cfg_is_fp16_d1[15] & (|in_dat_data_pack[254:250]);
    in_dat_norm[14] = cfg_is_fp16_d1[14] & (|in_dat_data_pack[238:234]);
    in_dat_norm[13] = cfg_is_fp16_d1[13] & (|in_dat_data_pack[222:218]);
    in_dat_norm[12] = cfg_is_fp16_d1[12] & (|in_dat_data_pack[206:202]);
    in_dat_norm[11] = cfg_is_fp16_d1[11] & (|in_dat_data_pack[190:186]);
    in_dat_norm[10] = cfg_is_fp16_d1[10] & (|in_dat_data_pack[174:170]);
    in_dat_norm[9] = cfg_is_fp16_d1[9] & (|in_dat_data_pack[158:154]);
    in_dat_norm[8] = cfg_is_fp16_d1[8] & (|in_dat_data_pack[142:138]);
    in_dat_norm[7] = cfg_is_fp16_d1[7] & (|in_dat_data_pack[126:122]);
    in_dat_norm[6] = cfg_is_fp16_d1[6] & (|in_dat_data_pack[110:106]);
    in_dat_norm[5] = cfg_is_fp16_d1[5] & (|in_dat_data_pack[94:90]);
    in_dat_norm[4] = cfg_is_fp16_d1[4] & (|in_dat_data_pack[78:74]);
    in_dat_norm[3] = cfg_is_fp16_d1[3] & (|in_dat_data_pack[62:58]);
    in_dat_norm[2] = cfg_is_fp16_d1[2] & (|in_dat_data_pack[46:42]);
    in_dat_norm[1] = cfg_is_fp16_d1[1] & (|in_dat_data_pack[30:26]);
    in_dat_norm[0] = cfg_is_fp16_d1[0] & (|in_dat_data_pack[14:10]);
end




always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori63 = ~cfg_is_fp16_d1[63] ? 12'b0 :
                                   in_dat_norm[63] ? {2'b1, in_dat_data_pack[1017:1008]} :
                                   {1'b0, in_dat_data_pack[1017:1008], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori62 = ~cfg_is_fp16_d1[62] ? 12'b0 :
                                   in_dat_norm[62] ? {2'b1, in_dat_data_pack[1001:992]} :
                                   {1'b0, in_dat_data_pack[1001:992], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori61 = ~cfg_is_fp16_d1[61] ? 12'b0 :
                                   in_dat_norm[61] ? {2'b1, in_dat_data_pack[985:976]} :
                                   {1'b0, in_dat_data_pack[985:976], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori60 = ~cfg_is_fp16_d1[60] ? 12'b0 :
                                   in_dat_norm[60] ? {2'b1, in_dat_data_pack[969:960]} :
                                   {1'b0, in_dat_data_pack[969:960], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori59 = ~cfg_is_fp16_d1[59] ? 12'b0 :
                                   in_dat_norm[59] ? {2'b1, in_dat_data_pack[953:944]} :
                                   {1'b0, in_dat_data_pack[953:944], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori58 = ~cfg_is_fp16_d1[58] ? 12'b0 :
                                   in_dat_norm[58] ? {2'b1, in_dat_data_pack[937:928]} :
                                   {1'b0, in_dat_data_pack[937:928], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori57 = ~cfg_is_fp16_d1[57] ? 12'b0 :
                                   in_dat_norm[57] ? {2'b1, in_dat_data_pack[921:912]} :
                                   {1'b0, in_dat_data_pack[921:912], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori56 = ~cfg_is_fp16_d1[56] ? 12'b0 :
                                   in_dat_norm[56] ? {2'b1, in_dat_data_pack[905:896]} :
                                   {1'b0, in_dat_data_pack[905:896], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori55 = ~cfg_is_fp16_d1[55] ? 12'b0 :
                                   in_dat_norm[55] ? {2'b1, in_dat_data_pack[889:880]} :
                                   {1'b0, in_dat_data_pack[889:880], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori54 = ~cfg_is_fp16_d1[54] ? 12'b0 :
                                   in_dat_norm[54] ? {2'b1, in_dat_data_pack[873:864]} :
                                   {1'b0, in_dat_data_pack[873:864], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori53 = ~cfg_is_fp16_d1[53] ? 12'b0 :
                                   in_dat_norm[53] ? {2'b1, in_dat_data_pack[857:848]} :
                                   {1'b0, in_dat_data_pack[857:848], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori52 = ~cfg_is_fp16_d1[52] ? 12'b0 :
                                   in_dat_norm[52] ? {2'b1, in_dat_data_pack[841:832]} :
                                   {1'b0, in_dat_data_pack[841:832], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori51 = ~cfg_is_fp16_d1[51] ? 12'b0 :
                                   in_dat_norm[51] ? {2'b1, in_dat_data_pack[825:816]} :
                                   {1'b0, in_dat_data_pack[825:816], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori50 = ~cfg_is_fp16_d1[50] ? 12'b0 :
                                   in_dat_norm[50] ? {2'b1, in_dat_data_pack[809:800]} :
                                   {1'b0, in_dat_data_pack[809:800], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori49 = ~cfg_is_fp16_d1[49] ? 12'b0 :
                                   in_dat_norm[49] ? {2'b1, in_dat_data_pack[793:784]} :
                                   {1'b0, in_dat_data_pack[793:784], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori48 = ~cfg_is_fp16_d1[48] ? 12'b0 :
                                   in_dat_norm[48] ? {2'b1, in_dat_data_pack[777:768]} :
                                   {1'b0, in_dat_data_pack[777:768], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori47 = ~cfg_is_fp16_d1[47] ? 12'b0 :
                                   in_dat_norm[47] ? {2'b1, in_dat_data_pack[761:752]} :
                                   {1'b0, in_dat_data_pack[761:752], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori46 = ~cfg_is_fp16_d1[46] ? 12'b0 :
                                   in_dat_norm[46] ? {2'b1, in_dat_data_pack[745:736]} :
                                   {1'b0, in_dat_data_pack[745:736], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori45 = ~cfg_is_fp16_d1[45] ? 12'b0 :
                                   in_dat_norm[45] ? {2'b1, in_dat_data_pack[729:720]} :
                                   {1'b0, in_dat_data_pack[729:720], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori44 = ~cfg_is_fp16_d1[44] ? 12'b0 :
                                   in_dat_norm[44] ? {2'b1, in_dat_data_pack[713:704]} :
                                   {1'b0, in_dat_data_pack[713:704], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori43 = ~cfg_is_fp16_d1[43] ? 12'b0 :
                                   in_dat_norm[43] ? {2'b1, in_dat_data_pack[697:688]} :
                                   {1'b0, in_dat_data_pack[697:688], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori42 = ~cfg_is_fp16_d1[42] ? 12'b0 :
                                   in_dat_norm[42] ? {2'b1, in_dat_data_pack[681:672]} :
                                   {1'b0, in_dat_data_pack[681:672], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori41 = ~cfg_is_fp16_d1[41] ? 12'b0 :
                                   in_dat_norm[41] ? {2'b1, in_dat_data_pack[665:656]} :
                                   {1'b0, in_dat_data_pack[665:656], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori40 = ~cfg_is_fp16_d1[40] ? 12'b0 :
                                   in_dat_norm[40] ? {2'b1, in_dat_data_pack[649:640]} :
                                   {1'b0, in_dat_data_pack[649:640], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori39 = ~cfg_is_fp16_d1[39] ? 12'b0 :
                                   in_dat_norm[39] ? {2'b1, in_dat_data_pack[633:624]} :
                                   {1'b0, in_dat_data_pack[633:624], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori38 = ~cfg_is_fp16_d1[38] ? 12'b0 :
                                   in_dat_norm[38] ? {2'b1, in_dat_data_pack[617:608]} :
                                   {1'b0, in_dat_data_pack[617:608], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori37 = ~cfg_is_fp16_d1[37] ? 12'b0 :
                                   in_dat_norm[37] ? {2'b1, in_dat_data_pack[601:592]} :
                                   {1'b0, in_dat_data_pack[601:592], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori36 = ~cfg_is_fp16_d1[36] ? 12'b0 :
                                   in_dat_norm[36] ? {2'b1, in_dat_data_pack[585:576]} :
                                   {1'b0, in_dat_data_pack[585:576], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori35 = ~cfg_is_fp16_d1[35] ? 12'b0 :
                                   in_dat_norm[35] ? {2'b1, in_dat_data_pack[569:560]} :
                                   {1'b0, in_dat_data_pack[569:560], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori34 = ~cfg_is_fp16_d1[34] ? 12'b0 :
                                   in_dat_norm[34] ? {2'b1, in_dat_data_pack[553:544]} :
                                   {1'b0, in_dat_data_pack[553:544], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori33 = ~cfg_is_fp16_d1[33] ? 12'b0 :
                                   in_dat_norm[33] ? {2'b1, in_dat_data_pack[537:528]} :
                                   {1'b0, in_dat_data_pack[537:528], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori32 = ~cfg_is_fp16_d1[32] ? 12'b0 :
                                   in_dat_norm[32] ? {2'b1, in_dat_data_pack[521:512]} :
                                   {1'b0, in_dat_data_pack[521:512], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori31 = ~cfg_is_fp16_d1[31] ? 12'b0 :
                                   in_dat_norm[31] ? {2'b1, in_dat_data_pack[505:496]} :
                                   {1'b0, in_dat_data_pack[505:496], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori30 = ~cfg_is_fp16_d1[30] ? 12'b0 :
                                   in_dat_norm[30] ? {2'b1, in_dat_data_pack[489:480]} :
                                   {1'b0, in_dat_data_pack[489:480], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori29 = ~cfg_is_fp16_d1[29] ? 12'b0 :
                                   in_dat_norm[29] ? {2'b1, in_dat_data_pack[473:464]} :
                                   {1'b0, in_dat_data_pack[473:464], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori28 = ~cfg_is_fp16_d1[28] ? 12'b0 :
                                   in_dat_norm[28] ? {2'b1, in_dat_data_pack[457:448]} :
                                   {1'b0, in_dat_data_pack[457:448], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori27 = ~cfg_is_fp16_d1[27] ? 12'b0 :
                                   in_dat_norm[27] ? {2'b1, in_dat_data_pack[441:432]} :
                                   {1'b0, in_dat_data_pack[441:432], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori26 = ~cfg_is_fp16_d1[26] ? 12'b0 :
                                   in_dat_norm[26] ? {2'b1, in_dat_data_pack[425:416]} :
                                   {1'b0, in_dat_data_pack[425:416], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori25 = ~cfg_is_fp16_d1[25] ? 12'b0 :
                                   in_dat_norm[25] ? {2'b1, in_dat_data_pack[409:400]} :
                                   {1'b0, in_dat_data_pack[409:400], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori24 = ~cfg_is_fp16_d1[24] ? 12'b0 :
                                   in_dat_norm[24] ? {2'b1, in_dat_data_pack[393:384]} :
                                   {1'b0, in_dat_data_pack[393:384], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori23 = ~cfg_is_fp16_d1[23] ? 12'b0 :
                                   in_dat_norm[23] ? {2'b1, in_dat_data_pack[377:368]} :
                                   {1'b0, in_dat_data_pack[377:368], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori22 = ~cfg_is_fp16_d1[22] ? 12'b0 :
                                   in_dat_norm[22] ? {2'b1, in_dat_data_pack[361:352]} :
                                   {1'b0, in_dat_data_pack[361:352], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori21 = ~cfg_is_fp16_d1[21] ? 12'b0 :
                                   in_dat_norm[21] ? {2'b1, in_dat_data_pack[345:336]} :
                                   {1'b0, in_dat_data_pack[345:336], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori20 = ~cfg_is_fp16_d1[20] ? 12'b0 :
                                   in_dat_norm[20] ? {2'b1, in_dat_data_pack[329:320]} :
                                   {1'b0, in_dat_data_pack[329:320], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori19 = ~cfg_is_fp16_d1[19] ? 12'b0 :
                                   in_dat_norm[19] ? {2'b1, in_dat_data_pack[313:304]} :
                                   {1'b0, in_dat_data_pack[313:304], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori18 = ~cfg_is_fp16_d1[18] ? 12'b0 :
                                   in_dat_norm[18] ? {2'b1, in_dat_data_pack[297:288]} :
                                   {1'b0, in_dat_data_pack[297:288], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori17 = ~cfg_is_fp16_d1[17] ? 12'b0 :
                                   in_dat_norm[17] ? {2'b1, in_dat_data_pack[281:272]} :
                                   {1'b0, in_dat_data_pack[281:272], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori16 = ~cfg_is_fp16_d1[16] ? 12'b0 :
                                   in_dat_norm[16] ? {2'b1, in_dat_data_pack[265:256]} :
                                   {1'b0, in_dat_data_pack[265:256], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori15 = ~cfg_is_fp16_d1[15] ? 12'b0 :
                                   in_dat_norm[15] ? {2'b1, in_dat_data_pack[249:240]} :
                                   {1'b0, in_dat_data_pack[249:240], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori14 = ~cfg_is_fp16_d1[14] ? 12'b0 :
                                   in_dat_norm[14] ? {2'b1, in_dat_data_pack[233:224]} :
                                   {1'b0, in_dat_data_pack[233:224], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori13 = ~cfg_is_fp16_d1[13] ? 12'b0 :
                                   in_dat_norm[13] ? {2'b1, in_dat_data_pack[217:208]} :
                                   {1'b0, in_dat_data_pack[217:208], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori12 = ~cfg_is_fp16_d1[12] ? 12'b0 :
                                   in_dat_norm[12] ? {2'b1, in_dat_data_pack[201:192]} :
                                   {1'b0, in_dat_data_pack[201:192], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori11 = ~cfg_is_fp16_d1[11] ? 12'b0 :
                                   in_dat_norm[11] ? {2'b1, in_dat_data_pack[185:176]} :
                                   {1'b0, in_dat_data_pack[185:176], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori10 = ~cfg_is_fp16_d1[10] ? 12'b0 :
                                   in_dat_norm[10] ? {2'b1, in_dat_data_pack[169:160]} :
                                   {1'b0, in_dat_data_pack[169:160], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori9 = ~cfg_is_fp16_d1[9] ? 12'b0 :
                                   in_dat_norm[9] ? {2'b1, in_dat_data_pack[153:144]} :
                                   {1'b0, in_dat_data_pack[153:144], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori8 = ~cfg_is_fp16_d1[8] ? 12'b0 :
                                   in_dat_norm[8] ? {2'b1, in_dat_data_pack[137:128]} :
                                   {1'b0, in_dat_data_pack[137:128], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori7 = ~cfg_is_fp16_d1[7] ? 12'b0 :
                                   in_dat_norm[7] ? {2'b1, in_dat_data_pack[121:112]} :
                                   {1'b0, in_dat_data_pack[121:112], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori6 = ~cfg_is_fp16_d1[6] ? 12'b0 :
                                   in_dat_norm[6] ? {2'b1, in_dat_data_pack[105:96]} :
                                   {1'b0, in_dat_data_pack[105:96], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori5 = ~cfg_is_fp16_d1[5] ? 12'b0 :
                                   in_dat_norm[5] ? {2'b1, in_dat_data_pack[89:80]} :
                                   {1'b0, in_dat_data_pack[89:80], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori4 = ~cfg_is_fp16_d1[4] ? 12'b0 :
                                   in_dat_norm[4] ? {2'b1, in_dat_data_pack[73:64]} :
                                   {1'b0, in_dat_data_pack[73:64], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori3 = ~cfg_is_fp16_d1[3] ? 12'b0 :
                                   in_dat_norm[3] ? {2'b1, in_dat_data_pack[57:48]} :
                                   {1'b0, in_dat_data_pack[57:48], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori2 = ~cfg_is_fp16_d1[2] ? 12'b0 :
                                   in_dat_norm[2] ? {2'b1, in_dat_data_pack[41:32]} :
                                   {1'b0, in_dat_data_pack[41:32], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori1 = ~cfg_is_fp16_d1[1] ? 12'b0 :
                                   in_dat_norm[1] ? {2'b1, in_dat_data_pack[25:16]} :
                                   {1'b0, in_dat_data_pack[25:16], 1'b0};
end



always @(
  cfg_is_fp16_d1
  or in_dat_norm
  or in_dat_data_pack
  ) begin
    in_dat_data_fp16_mts_ori0 = ~cfg_is_fp16_d1[0] ? 12'b0 :
                                   in_dat_norm[0] ? {2'b1, in_dat_data_pack[9:0]} :
                                   {1'b0, in_dat_data_pack[9:0], 1'b0};
end







always @(
  in_dat_data_fp16_mts_ori63
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft63[14:0] = ({3'b0, in_dat_data_fp16_mts_ori63} << in_dat_data_pack[1019:1018]);
    in_dat_data_fp16_63 = ({16{cfg_is_fp16_d1[63]}} & {in_dat_data_pack[1023], in_dat_data_fp16_mts_sft63});
end



always @(
  in_dat_data_fp16_mts_ori62
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft62[14:0] = ({3'b0, in_dat_data_fp16_mts_ori62} << in_dat_data_pack[1003:1002]);
    in_dat_data_fp16_62 = ({16{cfg_is_fp16_d1[62]}} & {in_dat_data_pack[1007], in_dat_data_fp16_mts_sft62});
end



always @(
  in_dat_data_fp16_mts_ori61
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft61[14:0] = ({3'b0, in_dat_data_fp16_mts_ori61} << in_dat_data_pack[987:986]);
    in_dat_data_fp16_61 = ({16{cfg_is_fp16_d1[61]}} & {in_dat_data_pack[991], in_dat_data_fp16_mts_sft61});
end



always @(
  in_dat_data_fp16_mts_ori60
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft60[14:0] = ({3'b0, in_dat_data_fp16_mts_ori60} << in_dat_data_pack[971:970]);
    in_dat_data_fp16_60 = ({16{cfg_is_fp16_d1[60]}} & {in_dat_data_pack[975], in_dat_data_fp16_mts_sft60});
end



always @(
  in_dat_data_fp16_mts_ori59
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft59[14:0] = ({3'b0, in_dat_data_fp16_mts_ori59} << in_dat_data_pack[955:954]);
    in_dat_data_fp16_59 = ({16{cfg_is_fp16_d1[59]}} & {in_dat_data_pack[959], in_dat_data_fp16_mts_sft59});
end



always @(
  in_dat_data_fp16_mts_ori58
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft58[14:0] = ({3'b0, in_dat_data_fp16_mts_ori58} << in_dat_data_pack[939:938]);
    in_dat_data_fp16_58 = ({16{cfg_is_fp16_d1[58]}} & {in_dat_data_pack[943], in_dat_data_fp16_mts_sft58});
end



always @(
  in_dat_data_fp16_mts_ori57
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft57[14:0] = ({3'b0, in_dat_data_fp16_mts_ori57} << in_dat_data_pack[923:922]);
    in_dat_data_fp16_57 = ({16{cfg_is_fp16_d1[57]}} & {in_dat_data_pack[927], in_dat_data_fp16_mts_sft57});
end



always @(
  in_dat_data_fp16_mts_ori56
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft56[14:0] = ({3'b0, in_dat_data_fp16_mts_ori56} << in_dat_data_pack[907:906]);
    in_dat_data_fp16_56 = ({16{cfg_is_fp16_d1[56]}} & {in_dat_data_pack[911], in_dat_data_fp16_mts_sft56});
end



always @(
  in_dat_data_fp16_mts_ori55
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft55[14:0] = ({3'b0, in_dat_data_fp16_mts_ori55} << in_dat_data_pack[891:890]);
    in_dat_data_fp16_55 = ({16{cfg_is_fp16_d1[55]}} & {in_dat_data_pack[895], in_dat_data_fp16_mts_sft55});
end



always @(
  in_dat_data_fp16_mts_ori54
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft54[14:0] = ({3'b0, in_dat_data_fp16_mts_ori54} << in_dat_data_pack[875:874]);
    in_dat_data_fp16_54 = ({16{cfg_is_fp16_d1[54]}} & {in_dat_data_pack[879], in_dat_data_fp16_mts_sft54});
end



always @(
  in_dat_data_fp16_mts_ori53
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft53[14:0] = ({3'b0, in_dat_data_fp16_mts_ori53} << in_dat_data_pack[859:858]);
    in_dat_data_fp16_53 = ({16{cfg_is_fp16_d1[53]}} & {in_dat_data_pack[863], in_dat_data_fp16_mts_sft53});
end



always @(
  in_dat_data_fp16_mts_ori52
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft52[14:0] = ({3'b0, in_dat_data_fp16_mts_ori52} << in_dat_data_pack[843:842]);
    in_dat_data_fp16_52 = ({16{cfg_is_fp16_d1[52]}} & {in_dat_data_pack[847], in_dat_data_fp16_mts_sft52});
end



always @(
  in_dat_data_fp16_mts_ori51
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft51[14:0] = ({3'b0, in_dat_data_fp16_mts_ori51} << in_dat_data_pack[827:826]);
    in_dat_data_fp16_51 = ({16{cfg_is_fp16_d1[51]}} & {in_dat_data_pack[831], in_dat_data_fp16_mts_sft51});
end



always @(
  in_dat_data_fp16_mts_ori50
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft50[14:0] = ({3'b0, in_dat_data_fp16_mts_ori50} << in_dat_data_pack[811:810]);
    in_dat_data_fp16_50 = ({16{cfg_is_fp16_d1[50]}} & {in_dat_data_pack[815], in_dat_data_fp16_mts_sft50});
end



always @(
  in_dat_data_fp16_mts_ori49
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft49[14:0] = ({3'b0, in_dat_data_fp16_mts_ori49} << in_dat_data_pack[795:794]);
    in_dat_data_fp16_49 = ({16{cfg_is_fp16_d1[49]}} & {in_dat_data_pack[799], in_dat_data_fp16_mts_sft49});
end



always @(
  in_dat_data_fp16_mts_ori48
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft48[14:0] = ({3'b0, in_dat_data_fp16_mts_ori48} << in_dat_data_pack[779:778]);
    in_dat_data_fp16_48 = ({16{cfg_is_fp16_d1[48]}} & {in_dat_data_pack[783], in_dat_data_fp16_mts_sft48});
end



always @(
  in_dat_data_fp16_mts_ori47
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft47[14:0] = ({3'b0, in_dat_data_fp16_mts_ori47} << in_dat_data_pack[763:762]);
    in_dat_data_fp16_47 = ({16{cfg_is_fp16_d1[47]}} & {in_dat_data_pack[767], in_dat_data_fp16_mts_sft47});
end



always @(
  in_dat_data_fp16_mts_ori46
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft46[14:0] = ({3'b0, in_dat_data_fp16_mts_ori46} << in_dat_data_pack[747:746]);
    in_dat_data_fp16_46 = ({16{cfg_is_fp16_d1[46]}} & {in_dat_data_pack[751], in_dat_data_fp16_mts_sft46});
end



always @(
  in_dat_data_fp16_mts_ori45
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft45[14:0] = ({3'b0, in_dat_data_fp16_mts_ori45} << in_dat_data_pack[731:730]);
    in_dat_data_fp16_45 = ({16{cfg_is_fp16_d1[45]}} & {in_dat_data_pack[735], in_dat_data_fp16_mts_sft45});
end



always @(
  in_dat_data_fp16_mts_ori44
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft44[14:0] = ({3'b0, in_dat_data_fp16_mts_ori44} << in_dat_data_pack[715:714]);
    in_dat_data_fp16_44 = ({16{cfg_is_fp16_d1[44]}} & {in_dat_data_pack[719], in_dat_data_fp16_mts_sft44});
end



always @(
  in_dat_data_fp16_mts_ori43
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft43[14:0] = ({3'b0, in_dat_data_fp16_mts_ori43} << in_dat_data_pack[699:698]);
    in_dat_data_fp16_43 = ({16{cfg_is_fp16_d1[43]}} & {in_dat_data_pack[703], in_dat_data_fp16_mts_sft43});
end



always @(
  in_dat_data_fp16_mts_ori42
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft42[14:0] = ({3'b0, in_dat_data_fp16_mts_ori42} << in_dat_data_pack[683:682]);
    in_dat_data_fp16_42 = ({16{cfg_is_fp16_d1[42]}} & {in_dat_data_pack[687], in_dat_data_fp16_mts_sft42});
end



always @(
  in_dat_data_fp16_mts_ori41
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft41[14:0] = ({3'b0, in_dat_data_fp16_mts_ori41} << in_dat_data_pack[667:666]);
    in_dat_data_fp16_41 = ({16{cfg_is_fp16_d1[41]}} & {in_dat_data_pack[671], in_dat_data_fp16_mts_sft41});
end



always @(
  in_dat_data_fp16_mts_ori40
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft40[14:0] = ({3'b0, in_dat_data_fp16_mts_ori40} << in_dat_data_pack[651:650]);
    in_dat_data_fp16_40 = ({16{cfg_is_fp16_d1[40]}} & {in_dat_data_pack[655], in_dat_data_fp16_mts_sft40});
end



always @(
  in_dat_data_fp16_mts_ori39
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft39[14:0] = ({3'b0, in_dat_data_fp16_mts_ori39} << in_dat_data_pack[635:634]);
    in_dat_data_fp16_39 = ({16{cfg_is_fp16_d1[39]}} & {in_dat_data_pack[639], in_dat_data_fp16_mts_sft39});
end



always @(
  in_dat_data_fp16_mts_ori38
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft38[14:0] = ({3'b0, in_dat_data_fp16_mts_ori38} << in_dat_data_pack[619:618]);
    in_dat_data_fp16_38 = ({16{cfg_is_fp16_d1[38]}} & {in_dat_data_pack[623], in_dat_data_fp16_mts_sft38});
end



always @(
  in_dat_data_fp16_mts_ori37
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft37[14:0] = ({3'b0, in_dat_data_fp16_mts_ori37} << in_dat_data_pack[603:602]);
    in_dat_data_fp16_37 = ({16{cfg_is_fp16_d1[37]}} & {in_dat_data_pack[607], in_dat_data_fp16_mts_sft37});
end



always @(
  in_dat_data_fp16_mts_ori36
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft36[14:0] = ({3'b0, in_dat_data_fp16_mts_ori36} << in_dat_data_pack[587:586]);
    in_dat_data_fp16_36 = ({16{cfg_is_fp16_d1[36]}} & {in_dat_data_pack[591], in_dat_data_fp16_mts_sft36});
end



always @(
  in_dat_data_fp16_mts_ori35
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft35[14:0] = ({3'b0, in_dat_data_fp16_mts_ori35} << in_dat_data_pack[571:570]);
    in_dat_data_fp16_35 = ({16{cfg_is_fp16_d1[35]}} & {in_dat_data_pack[575], in_dat_data_fp16_mts_sft35});
end



always @(
  in_dat_data_fp16_mts_ori34
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft34[14:0] = ({3'b0, in_dat_data_fp16_mts_ori34} << in_dat_data_pack[555:554]);
    in_dat_data_fp16_34 = ({16{cfg_is_fp16_d1[34]}} & {in_dat_data_pack[559], in_dat_data_fp16_mts_sft34});
end



always @(
  in_dat_data_fp16_mts_ori33
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft33[14:0] = ({3'b0, in_dat_data_fp16_mts_ori33} << in_dat_data_pack[539:538]);
    in_dat_data_fp16_33 = ({16{cfg_is_fp16_d1[33]}} & {in_dat_data_pack[543], in_dat_data_fp16_mts_sft33});
end



always @(
  in_dat_data_fp16_mts_ori32
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft32[14:0] = ({3'b0, in_dat_data_fp16_mts_ori32} << in_dat_data_pack[523:522]);
    in_dat_data_fp16_32 = ({16{cfg_is_fp16_d1[32]}} & {in_dat_data_pack[527], in_dat_data_fp16_mts_sft32});
end



always @(
  in_dat_data_fp16_mts_ori31
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft31[14:0] = ({3'b0, in_dat_data_fp16_mts_ori31} << in_dat_data_pack[507:506]);
    in_dat_data_fp16_31 = ({16{cfg_is_fp16_d1[31]}} & {in_dat_data_pack[511], in_dat_data_fp16_mts_sft31});
end



always @(
  in_dat_data_fp16_mts_ori30
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft30[14:0] = ({3'b0, in_dat_data_fp16_mts_ori30} << in_dat_data_pack[491:490]);
    in_dat_data_fp16_30 = ({16{cfg_is_fp16_d1[30]}} & {in_dat_data_pack[495], in_dat_data_fp16_mts_sft30});
end



always @(
  in_dat_data_fp16_mts_ori29
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft29[14:0] = ({3'b0, in_dat_data_fp16_mts_ori29} << in_dat_data_pack[475:474]);
    in_dat_data_fp16_29 = ({16{cfg_is_fp16_d1[29]}} & {in_dat_data_pack[479], in_dat_data_fp16_mts_sft29});
end



always @(
  in_dat_data_fp16_mts_ori28
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft28[14:0] = ({3'b0, in_dat_data_fp16_mts_ori28} << in_dat_data_pack[459:458]);
    in_dat_data_fp16_28 = ({16{cfg_is_fp16_d1[28]}} & {in_dat_data_pack[463], in_dat_data_fp16_mts_sft28});
end



always @(
  in_dat_data_fp16_mts_ori27
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft27[14:0] = ({3'b0, in_dat_data_fp16_mts_ori27} << in_dat_data_pack[443:442]);
    in_dat_data_fp16_27 = ({16{cfg_is_fp16_d1[27]}} & {in_dat_data_pack[447], in_dat_data_fp16_mts_sft27});
end



always @(
  in_dat_data_fp16_mts_ori26
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft26[14:0] = ({3'b0, in_dat_data_fp16_mts_ori26} << in_dat_data_pack[427:426]);
    in_dat_data_fp16_26 = ({16{cfg_is_fp16_d1[26]}} & {in_dat_data_pack[431], in_dat_data_fp16_mts_sft26});
end



always @(
  in_dat_data_fp16_mts_ori25
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft25[14:0] = ({3'b0, in_dat_data_fp16_mts_ori25} << in_dat_data_pack[411:410]);
    in_dat_data_fp16_25 = ({16{cfg_is_fp16_d1[25]}} & {in_dat_data_pack[415], in_dat_data_fp16_mts_sft25});
end



always @(
  in_dat_data_fp16_mts_ori24
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft24[14:0] = ({3'b0, in_dat_data_fp16_mts_ori24} << in_dat_data_pack[395:394]);
    in_dat_data_fp16_24 = ({16{cfg_is_fp16_d1[24]}} & {in_dat_data_pack[399], in_dat_data_fp16_mts_sft24});
end



always @(
  in_dat_data_fp16_mts_ori23
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft23[14:0] = ({3'b0, in_dat_data_fp16_mts_ori23} << in_dat_data_pack[379:378]);
    in_dat_data_fp16_23 = ({16{cfg_is_fp16_d1[23]}} & {in_dat_data_pack[383], in_dat_data_fp16_mts_sft23});
end



always @(
  in_dat_data_fp16_mts_ori22
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft22[14:0] = ({3'b0, in_dat_data_fp16_mts_ori22} << in_dat_data_pack[363:362]);
    in_dat_data_fp16_22 = ({16{cfg_is_fp16_d1[22]}} & {in_dat_data_pack[367], in_dat_data_fp16_mts_sft22});
end



always @(
  in_dat_data_fp16_mts_ori21
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft21[14:0] = ({3'b0, in_dat_data_fp16_mts_ori21} << in_dat_data_pack[347:346]);
    in_dat_data_fp16_21 = ({16{cfg_is_fp16_d1[21]}} & {in_dat_data_pack[351], in_dat_data_fp16_mts_sft21});
end



always @(
  in_dat_data_fp16_mts_ori20
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft20[14:0] = ({3'b0, in_dat_data_fp16_mts_ori20} << in_dat_data_pack[331:330]);
    in_dat_data_fp16_20 = ({16{cfg_is_fp16_d1[20]}} & {in_dat_data_pack[335], in_dat_data_fp16_mts_sft20});
end



always @(
  in_dat_data_fp16_mts_ori19
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft19[14:0] = ({3'b0, in_dat_data_fp16_mts_ori19} << in_dat_data_pack[315:314]);
    in_dat_data_fp16_19 = ({16{cfg_is_fp16_d1[19]}} & {in_dat_data_pack[319], in_dat_data_fp16_mts_sft19});
end



always @(
  in_dat_data_fp16_mts_ori18
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft18[14:0] = ({3'b0, in_dat_data_fp16_mts_ori18} << in_dat_data_pack[299:298]);
    in_dat_data_fp16_18 = ({16{cfg_is_fp16_d1[18]}} & {in_dat_data_pack[303], in_dat_data_fp16_mts_sft18});
end



always @(
  in_dat_data_fp16_mts_ori17
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft17[14:0] = ({3'b0, in_dat_data_fp16_mts_ori17} << in_dat_data_pack[283:282]);
    in_dat_data_fp16_17 = ({16{cfg_is_fp16_d1[17]}} & {in_dat_data_pack[287], in_dat_data_fp16_mts_sft17});
end



always @(
  in_dat_data_fp16_mts_ori16
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft16[14:0] = ({3'b0, in_dat_data_fp16_mts_ori16} << in_dat_data_pack[267:266]);
    in_dat_data_fp16_16 = ({16{cfg_is_fp16_d1[16]}} & {in_dat_data_pack[271], in_dat_data_fp16_mts_sft16});
end



always @(
  in_dat_data_fp16_mts_ori15
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft15[14:0] = ({3'b0, in_dat_data_fp16_mts_ori15} << in_dat_data_pack[251:250]);
    in_dat_data_fp16_15 = ({16{cfg_is_fp16_d1[15]}} & {in_dat_data_pack[255], in_dat_data_fp16_mts_sft15});
end



always @(
  in_dat_data_fp16_mts_ori14
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft14[14:0] = ({3'b0, in_dat_data_fp16_mts_ori14} << in_dat_data_pack[235:234]);
    in_dat_data_fp16_14 = ({16{cfg_is_fp16_d1[14]}} & {in_dat_data_pack[239], in_dat_data_fp16_mts_sft14});
end



always @(
  in_dat_data_fp16_mts_ori13
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft13[14:0] = ({3'b0, in_dat_data_fp16_mts_ori13} << in_dat_data_pack[219:218]);
    in_dat_data_fp16_13 = ({16{cfg_is_fp16_d1[13]}} & {in_dat_data_pack[223], in_dat_data_fp16_mts_sft13});
end



always @(
  in_dat_data_fp16_mts_ori12
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft12[14:0] = ({3'b0, in_dat_data_fp16_mts_ori12} << in_dat_data_pack[203:202]);
    in_dat_data_fp16_12 = ({16{cfg_is_fp16_d1[12]}} & {in_dat_data_pack[207], in_dat_data_fp16_mts_sft12});
end



always @(
  in_dat_data_fp16_mts_ori11
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft11[14:0] = ({3'b0, in_dat_data_fp16_mts_ori11} << in_dat_data_pack[187:186]);
    in_dat_data_fp16_11 = ({16{cfg_is_fp16_d1[11]}} & {in_dat_data_pack[191], in_dat_data_fp16_mts_sft11});
end



always @(
  in_dat_data_fp16_mts_ori10
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft10[14:0] = ({3'b0, in_dat_data_fp16_mts_ori10} << in_dat_data_pack[171:170]);
    in_dat_data_fp16_10 = ({16{cfg_is_fp16_d1[10]}} & {in_dat_data_pack[175], in_dat_data_fp16_mts_sft10});
end



always @(
  in_dat_data_fp16_mts_ori9
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft9[14:0] = ({3'b0, in_dat_data_fp16_mts_ori9} << in_dat_data_pack[155:154]);
    in_dat_data_fp16_9 = ({16{cfg_is_fp16_d1[9]}} & {in_dat_data_pack[159], in_dat_data_fp16_mts_sft9});
end



always @(
  in_dat_data_fp16_mts_ori8
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft8[14:0] = ({3'b0, in_dat_data_fp16_mts_ori8} << in_dat_data_pack[139:138]);
    in_dat_data_fp16_8 = ({16{cfg_is_fp16_d1[8]}} & {in_dat_data_pack[143], in_dat_data_fp16_mts_sft8});
end



always @(
  in_dat_data_fp16_mts_ori7
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft7[14:0] = ({3'b0, in_dat_data_fp16_mts_ori7} << in_dat_data_pack[123:122]);
    in_dat_data_fp16_7 = ({16{cfg_is_fp16_d1[7]}} & {in_dat_data_pack[127], in_dat_data_fp16_mts_sft7});
end



always @(
  in_dat_data_fp16_mts_ori6
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft6[14:0] = ({3'b0, in_dat_data_fp16_mts_ori6} << in_dat_data_pack[107:106]);
    in_dat_data_fp16_6 = ({16{cfg_is_fp16_d1[6]}} & {in_dat_data_pack[111], in_dat_data_fp16_mts_sft6});
end



always @(
  in_dat_data_fp16_mts_ori5
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft5[14:0] = ({3'b0, in_dat_data_fp16_mts_ori5} << in_dat_data_pack[91:90]);
    in_dat_data_fp16_5 = ({16{cfg_is_fp16_d1[5]}} & {in_dat_data_pack[95], in_dat_data_fp16_mts_sft5});
end



always @(
  in_dat_data_fp16_mts_ori4
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft4[14:0] = ({3'b0, in_dat_data_fp16_mts_ori4} << in_dat_data_pack[75:74]);
    in_dat_data_fp16_4 = ({16{cfg_is_fp16_d1[4]}} & {in_dat_data_pack[79], in_dat_data_fp16_mts_sft4});
end



always @(
  in_dat_data_fp16_mts_ori3
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft3[14:0] = ({3'b0, in_dat_data_fp16_mts_ori3} << in_dat_data_pack[59:58]);
    in_dat_data_fp16_3 = ({16{cfg_is_fp16_d1[3]}} & {in_dat_data_pack[63], in_dat_data_fp16_mts_sft3});
end



always @(
  in_dat_data_fp16_mts_ori2
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft2[14:0] = ({3'b0, in_dat_data_fp16_mts_ori2} << in_dat_data_pack[43:42]);
    in_dat_data_fp16_2 = ({16{cfg_is_fp16_d1[2]}} & {in_dat_data_pack[47], in_dat_data_fp16_mts_sft2});
end



always @(
  in_dat_data_fp16_mts_ori1
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft1[14:0] = ({3'b0, in_dat_data_fp16_mts_ori1} << in_dat_data_pack[27:26]);
    in_dat_data_fp16_1 = ({16{cfg_is_fp16_d1[1]}} & {in_dat_data_pack[31], in_dat_data_fp16_mts_sft1});
end



always @(
  in_dat_data_fp16_mts_ori0
  or in_dat_data_pack
  or cfg_is_fp16_d1
  ) begin
    in_dat_data_fp16_mts_sft0[14:0] = ({3'b0, in_dat_data_fp16_mts_ori0} << in_dat_data_pack[11:10]);
    in_dat_data_fp16_0 = ({16{cfg_is_fp16_d1[0]}} & {in_dat_data_pack[15], in_dat_data_fp16_mts_sft0});
end







always @(
  in_dat_nan
  ) begin
    dat_has_nan = (|in_dat_nan);
end

always @(
  in_dat_data_fp16_63
  or in_dat_data_fp16_62
  or in_dat_data_fp16_61
  or in_dat_data_fp16_60
  or in_dat_data_fp16_59
  or in_dat_data_fp16_58
  or in_dat_data_fp16_57
  or in_dat_data_fp16_56
  or in_dat_data_fp16_55
  or in_dat_data_fp16_54
  or in_dat_data_fp16_53
  or in_dat_data_fp16_52
  or in_dat_data_fp16_51
  or in_dat_data_fp16_50
  or in_dat_data_fp16_49
  or in_dat_data_fp16_48
  or in_dat_data_fp16_47
  or in_dat_data_fp16_46
  or in_dat_data_fp16_45
  or in_dat_data_fp16_44
  or in_dat_data_fp16_43
  or in_dat_data_fp16_42
  or in_dat_data_fp16_41
  or in_dat_data_fp16_40
  or in_dat_data_fp16_39
  or in_dat_data_fp16_38
  or in_dat_data_fp16_37
  or in_dat_data_fp16_36
  or in_dat_data_fp16_35
  or in_dat_data_fp16_34
  or in_dat_data_fp16_33
  or in_dat_data_fp16_32
  or in_dat_data_fp16_31
  or in_dat_data_fp16_30
  or in_dat_data_fp16_29
  or in_dat_data_fp16_28
  or in_dat_data_fp16_27
  or in_dat_data_fp16_26
  or in_dat_data_fp16_25
  or in_dat_data_fp16_24
  or in_dat_data_fp16_23
  or in_dat_data_fp16_22
  or in_dat_data_fp16_21
  or in_dat_data_fp16_20
  or in_dat_data_fp16_19
  or in_dat_data_fp16_18
  or in_dat_data_fp16_17
  or in_dat_data_fp16_16
  or in_dat_data_fp16_15
  or in_dat_data_fp16_14
  or in_dat_data_fp16_13
  or in_dat_data_fp16_12
  or in_dat_data_fp16_11
  or in_dat_data_fp16_10
  or in_dat_data_fp16_9
  or in_dat_data_fp16_8
  or in_dat_data_fp16_7
  or in_dat_data_fp16_6
  or in_dat_data_fp16_5
  or in_dat_data_fp16_4
  or in_dat_data_fp16_3
  or in_dat_data_fp16_2
  or in_dat_data_fp16_1
  or in_dat_data_fp16_0
  ) begin
    in_dat_data_fp16 = {in_dat_data_fp16_63, in_dat_data_fp16_62, in_dat_data_fp16_61, in_dat_data_fp16_60, in_dat_data_fp16_59, in_dat_data_fp16_58, in_dat_data_fp16_57, in_dat_data_fp16_56, in_dat_data_fp16_55, in_dat_data_fp16_54, in_dat_data_fp16_53, in_dat_data_fp16_52, in_dat_data_fp16_51, in_dat_data_fp16_50, in_dat_data_fp16_49, in_dat_data_fp16_48, in_dat_data_fp16_47, in_dat_data_fp16_46, in_dat_data_fp16_45, in_dat_data_fp16_44, in_dat_data_fp16_43, in_dat_data_fp16_42, in_dat_data_fp16_41, in_dat_data_fp16_40, in_dat_data_fp16_39, in_dat_data_fp16_38, in_dat_data_fp16_37, in_dat_data_fp16_36, in_dat_data_fp16_35, in_dat_data_fp16_34, in_dat_data_fp16_33, in_dat_data_fp16_32, in_dat_data_fp16_31, in_dat_data_fp16_30, in_dat_data_fp16_29, in_dat_data_fp16_28, in_dat_data_fp16_27, in_dat_data_fp16_26, in_dat_data_fp16_25, in_dat_data_fp16_24, in_dat_data_fp16_23, in_dat_data_fp16_22, in_dat_data_fp16_21, in_dat_data_fp16_20, in_dat_data_fp16_19, in_dat_data_fp16_18, in_dat_data_fp16_17, in_dat_data_fp16_16, in_dat_data_fp16_15, in_dat_data_fp16_14, in_dat_data_fp16_13, in_dat_data_fp16_12, in_dat_data_fp16_11, in_dat_data_fp16_10, in_dat_data_fp16_9, in_dat_data_fp16_8, in_dat_data_fp16_7, in_dat_data_fp16_6, in_dat_data_fp16_5, in_dat_data_fp16_4, in_dat_data_fp16_3, in_dat_data_fp16_2, in_dat_data_fp16_1, in_dat_data_fp16_0};
end

//////////////// dat_pre_data_w ////////////////
always @(
  in_dat_data_fp16
  or in_dat_data_int8
  or in_dat_data_int16
  ) begin
    dat_pre_data_w = in_dat_data_fp16 | in_dat_data_int8 | in_dat_data_int16;
end

always @(
  cfg_is_fp16_d1
  or dat_has_nan
  or in_dat_mask
  or cfg_is_int8_d1
  or in_dat_mask_int8
  ) begin
    dat_pre_nz_w = (cfg_is_fp16_d1[64]) ? {128{~dat_has_nan}} & in_dat_mask :
                   (cfg_is_int8_d1[64]) ? in_dat_mask_int8 :
                   in_dat_mask;
end

always @(
  in_dat_exp
  ) begin
    dat_pre_exp_w = in_dat_exp;
end

always @(
  dat_pre_nz_w
  ) begin
    dat_pre_mask_w = {dat_pre_nz_w[63*2],dat_pre_nz_w[62*2],dat_pre_nz_w[61*2],dat_pre_nz_w[60*2],dat_pre_nz_w[59*2],dat_pre_nz_w[58*2],dat_pre_nz_w[57*2],dat_pre_nz_w[56*2],dat_pre_nz_w[55*2],dat_pre_nz_w[54*2],dat_pre_nz_w[53*2],dat_pre_nz_w[52*2],dat_pre_nz_w[51*2],dat_pre_nz_w[50*2],dat_pre_nz_w[49*2],dat_pre_nz_w[48*2],dat_pre_nz_w[47*2],dat_pre_nz_w[46*2],dat_pre_nz_w[45*2],dat_pre_nz_w[44*2],dat_pre_nz_w[43*2],dat_pre_nz_w[42*2],dat_pre_nz_w[41*2],dat_pre_nz_w[40*2],dat_pre_nz_w[39*2],dat_pre_nz_w[38*2],dat_pre_nz_w[37*2],dat_pre_nz_w[36*2],dat_pre_nz_w[35*2],dat_pre_nz_w[34*2],dat_pre_nz_w[33*2],dat_pre_nz_w[32*2],dat_pre_nz_w[31*2],dat_pre_nz_w[30*2],dat_pre_nz_w[29*2],dat_pre_nz_w[28*2],dat_pre_nz_w[27*2],dat_pre_nz_w[26*2],dat_pre_nz_w[25*2],dat_pre_nz_w[24*2],dat_pre_nz_w[23*2],dat_pre_nz_w[22*2],dat_pre_nz_w[21*2],dat_pre_nz_w[20*2],dat_pre_nz_w[19*2],dat_pre_nz_w[18*2],dat_pre_nz_w[17*2],dat_pre_nz_w[16*2],dat_pre_nz_w[15*2],dat_pre_nz_w[14*2],dat_pre_nz_w[13*2],dat_pre_nz_w[12*2],dat_pre_nz_w[11*2],dat_pre_nz_w[10*2],dat_pre_nz_w[9*2],dat_pre_nz_w[8*2],dat_pre_nz_w[7*2],dat_pre_nz_w[6*2],dat_pre_nz_w[5*2],dat_pre_nz_w[4*2],dat_pre_nz_w[3*2],dat_pre_nz_w[2*2],dat_pre_nz_w[1*2],dat_pre_nz_w[0*2]};
end

//==========================================================
// Data pre-process register         
//==========================================================
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_pre_pvld <= {16{1'b0}};
  end else begin
  dat_pre_pvld <= {16{in_dat_pvld}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld) == 1'b1) begin
    dat_pre_nz <= dat_pre_nz_w;
  // VCS coverage off
  end else if ((in_dat_pvld) == 1'b0) begin
  end else begin
    dat_pre_nz <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[65]) == 1'b1) begin
    dat_pre_nan <= in_dat_nan;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[65]) == 1'b0) begin
  end else begin
    dat_pre_nan <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[0] | in_dat_nan[0])) == 1'b1) begin
    dat_pre_data[7:0] <= dat_pre_data_w[7:0];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[0] | in_dat_nan[0])) == 1'b0) begin
  end else begin
    dat_pre_data[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[1] | in_dat_nan[0])) == 1'b1) begin
    dat_pre_data[15:8] <= dat_pre_data_w[15:8];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[1] | in_dat_nan[0])) == 1'b0) begin
  end else begin
    dat_pre_data[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[2] | in_dat_nan[1])) == 1'b1) begin
    dat_pre_data[23:16] <= dat_pre_data_w[23:16];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[2] | in_dat_nan[1])) == 1'b0) begin
  end else begin
    dat_pre_data[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[3] | in_dat_nan[1])) == 1'b1) begin
    dat_pre_data[31:24] <= dat_pre_data_w[31:24];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[3] | in_dat_nan[1])) == 1'b0) begin
  end else begin
    dat_pre_data[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[4] | in_dat_nan[2])) == 1'b1) begin
    dat_pre_data[39:32] <= dat_pre_data_w[39:32];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[4] | in_dat_nan[2])) == 1'b0) begin
  end else begin
    dat_pre_data[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[5] | in_dat_nan[2])) == 1'b1) begin
    dat_pre_data[47:40] <= dat_pre_data_w[47:40];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[5] | in_dat_nan[2])) == 1'b0) begin
  end else begin
    dat_pre_data[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[6] | in_dat_nan[3])) == 1'b1) begin
    dat_pre_data[55:48] <= dat_pre_data_w[55:48];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[6] | in_dat_nan[3])) == 1'b0) begin
  end else begin
    dat_pre_data[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[7] | in_dat_nan[3])) == 1'b1) begin
    dat_pre_data[63:56] <= dat_pre_data_w[63:56];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[7] | in_dat_nan[3])) == 1'b0) begin
  end else begin
    dat_pre_data[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[8] | in_dat_nan[4])) == 1'b1) begin
    dat_pre_data[71:64] <= dat_pre_data_w[71:64];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[8] | in_dat_nan[4])) == 1'b0) begin
  end else begin
    dat_pre_data[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[9] | in_dat_nan[4])) == 1'b1) begin
    dat_pre_data[79:72] <= dat_pre_data_w[79:72];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[9] | in_dat_nan[4])) == 1'b0) begin
  end else begin
    dat_pre_data[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[10] | in_dat_nan[5])) == 1'b1) begin
    dat_pre_data[87:80] <= dat_pre_data_w[87:80];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[10] | in_dat_nan[5])) == 1'b0) begin
  end else begin
    dat_pre_data[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[11] | in_dat_nan[5])) == 1'b1) begin
    dat_pre_data[95:88] <= dat_pre_data_w[95:88];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[11] | in_dat_nan[5])) == 1'b0) begin
  end else begin
    dat_pre_data[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[12] | in_dat_nan[6])) == 1'b1) begin
    dat_pre_data[103:96] <= dat_pre_data_w[103:96];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[12] | in_dat_nan[6])) == 1'b0) begin
  end else begin
    dat_pre_data[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[13] | in_dat_nan[6])) == 1'b1) begin
    dat_pre_data[111:104] <= dat_pre_data_w[111:104];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[13] | in_dat_nan[6])) == 1'b0) begin
  end else begin
    dat_pre_data[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[14] | in_dat_nan[7])) == 1'b1) begin
    dat_pre_data[119:112] <= dat_pre_data_w[119:112];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[14] | in_dat_nan[7])) == 1'b0) begin
  end else begin
    dat_pre_data[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[15] | in_dat_nan[7])) == 1'b1) begin
    dat_pre_data[127:120] <= dat_pre_data_w[127:120];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[15] | in_dat_nan[7])) == 1'b0) begin
  end else begin
    dat_pre_data[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[16] | in_dat_nan[8])) == 1'b1) begin
    dat_pre_data[135:128] <= dat_pre_data_w[135:128];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[16] | in_dat_nan[8])) == 1'b0) begin
  end else begin
    dat_pre_data[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[17] | in_dat_nan[8])) == 1'b1) begin
    dat_pre_data[143:136] <= dat_pre_data_w[143:136];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[17] | in_dat_nan[8])) == 1'b0) begin
  end else begin
    dat_pre_data[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[18] | in_dat_nan[9])) == 1'b1) begin
    dat_pre_data[151:144] <= dat_pre_data_w[151:144];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[18] | in_dat_nan[9])) == 1'b0) begin
  end else begin
    dat_pre_data[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[19] | in_dat_nan[9])) == 1'b1) begin
    dat_pre_data[159:152] <= dat_pre_data_w[159:152];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[19] | in_dat_nan[9])) == 1'b0) begin
  end else begin
    dat_pre_data[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[20] | in_dat_nan[10])) == 1'b1) begin
    dat_pre_data[167:160] <= dat_pre_data_w[167:160];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[20] | in_dat_nan[10])) == 1'b0) begin
  end else begin
    dat_pre_data[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[21] | in_dat_nan[10])) == 1'b1) begin
    dat_pre_data[175:168] <= dat_pre_data_w[175:168];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[21] | in_dat_nan[10])) == 1'b0) begin
  end else begin
    dat_pre_data[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[22] | in_dat_nan[11])) == 1'b1) begin
    dat_pre_data[183:176] <= dat_pre_data_w[183:176];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[22] | in_dat_nan[11])) == 1'b0) begin
  end else begin
    dat_pre_data[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[23] | in_dat_nan[11])) == 1'b1) begin
    dat_pre_data[191:184] <= dat_pre_data_w[191:184];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[23] | in_dat_nan[11])) == 1'b0) begin
  end else begin
    dat_pre_data[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[24] | in_dat_nan[12])) == 1'b1) begin
    dat_pre_data[199:192] <= dat_pre_data_w[199:192];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[24] | in_dat_nan[12])) == 1'b0) begin
  end else begin
    dat_pre_data[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[25] | in_dat_nan[12])) == 1'b1) begin
    dat_pre_data[207:200] <= dat_pre_data_w[207:200];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[25] | in_dat_nan[12])) == 1'b0) begin
  end else begin
    dat_pre_data[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[26] | in_dat_nan[13])) == 1'b1) begin
    dat_pre_data[215:208] <= dat_pre_data_w[215:208];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[26] | in_dat_nan[13])) == 1'b0) begin
  end else begin
    dat_pre_data[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[27] | in_dat_nan[13])) == 1'b1) begin
    dat_pre_data[223:216] <= dat_pre_data_w[223:216];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[27] | in_dat_nan[13])) == 1'b0) begin
  end else begin
    dat_pre_data[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[28] | in_dat_nan[14])) == 1'b1) begin
    dat_pre_data[231:224] <= dat_pre_data_w[231:224];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[28] | in_dat_nan[14])) == 1'b0) begin
  end else begin
    dat_pre_data[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[29] | in_dat_nan[14])) == 1'b1) begin
    dat_pre_data[239:232] <= dat_pre_data_w[239:232];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[29] | in_dat_nan[14])) == 1'b0) begin
  end else begin
    dat_pre_data[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[30] | in_dat_nan[15])) == 1'b1) begin
    dat_pre_data[247:240] <= dat_pre_data_w[247:240];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[30] | in_dat_nan[15])) == 1'b0) begin
  end else begin
    dat_pre_data[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[31] | in_dat_nan[15])) == 1'b1) begin
    dat_pre_data[255:248] <= dat_pre_data_w[255:248];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[31] | in_dat_nan[15])) == 1'b0) begin
  end else begin
    dat_pre_data[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[32] | in_dat_nan[16])) == 1'b1) begin
    dat_pre_data[263:256] <= dat_pre_data_w[263:256];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[32] | in_dat_nan[16])) == 1'b0) begin
  end else begin
    dat_pre_data[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[33] | in_dat_nan[16])) == 1'b1) begin
    dat_pre_data[271:264] <= dat_pre_data_w[271:264];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[33] | in_dat_nan[16])) == 1'b0) begin
  end else begin
    dat_pre_data[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[34] | in_dat_nan[17])) == 1'b1) begin
    dat_pre_data[279:272] <= dat_pre_data_w[279:272];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[34] | in_dat_nan[17])) == 1'b0) begin
  end else begin
    dat_pre_data[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[35] | in_dat_nan[17])) == 1'b1) begin
    dat_pre_data[287:280] <= dat_pre_data_w[287:280];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[35] | in_dat_nan[17])) == 1'b0) begin
  end else begin
    dat_pre_data[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[36] | in_dat_nan[18])) == 1'b1) begin
    dat_pre_data[295:288] <= dat_pre_data_w[295:288];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[36] | in_dat_nan[18])) == 1'b0) begin
  end else begin
    dat_pre_data[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[37] | in_dat_nan[18])) == 1'b1) begin
    dat_pre_data[303:296] <= dat_pre_data_w[303:296];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[37] | in_dat_nan[18])) == 1'b0) begin
  end else begin
    dat_pre_data[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[38] | in_dat_nan[19])) == 1'b1) begin
    dat_pre_data[311:304] <= dat_pre_data_w[311:304];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[38] | in_dat_nan[19])) == 1'b0) begin
  end else begin
    dat_pre_data[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[39] | in_dat_nan[19])) == 1'b1) begin
    dat_pre_data[319:312] <= dat_pre_data_w[319:312];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[39] | in_dat_nan[19])) == 1'b0) begin
  end else begin
    dat_pre_data[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[40] | in_dat_nan[20])) == 1'b1) begin
    dat_pre_data[327:320] <= dat_pre_data_w[327:320];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[40] | in_dat_nan[20])) == 1'b0) begin
  end else begin
    dat_pre_data[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[41] | in_dat_nan[20])) == 1'b1) begin
    dat_pre_data[335:328] <= dat_pre_data_w[335:328];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[41] | in_dat_nan[20])) == 1'b0) begin
  end else begin
    dat_pre_data[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[42] | in_dat_nan[21])) == 1'b1) begin
    dat_pre_data[343:336] <= dat_pre_data_w[343:336];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[42] | in_dat_nan[21])) == 1'b0) begin
  end else begin
    dat_pre_data[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[43] | in_dat_nan[21])) == 1'b1) begin
    dat_pre_data[351:344] <= dat_pre_data_w[351:344];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[43] | in_dat_nan[21])) == 1'b0) begin
  end else begin
    dat_pre_data[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[44] | in_dat_nan[22])) == 1'b1) begin
    dat_pre_data[359:352] <= dat_pre_data_w[359:352];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[44] | in_dat_nan[22])) == 1'b0) begin
  end else begin
    dat_pre_data[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[45] | in_dat_nan[22])) == 1'b1) begin
    dat_pre_data[367:360] <= dat_pre_data_w[367:360];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[45] | in_dat_nan[22])) == 1'b0) begin
  end else begin
    dat_pre_data[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[46] | in_dat_nan[23])) == 1'b1) begin
    dat_pre_data[375:368] <= dat_pre_data_w[375:368];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[46] | in_dat_nan[23])) == 1'b0) begin
  end else begin
    dat_pre_data[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[47] | in_dat_nan[23])) == 1'b1) begin
    dat_pre_data[383:376] <= dat_pre_data_w[383:376];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[47] | in_dat_nan[23])) == 1'b0) begin
  end else begin
    dat_pre_data[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[48] | in_dat_nan[24])) == 1'b1) begin
    dat_pre_data[391:384] <= dat_pre_data_w[391:384];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[48] | in_dat_nan[24])) == 1'b0) begin
  end else begin
    dat_pre_data[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[49] | in_dat_nan[24])) == 1'b1) begin
    dat_pre_data[399:392] <= dat_pre_data_w[399:392];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[49] | in_dat_nan[24])) == 1'b0) begin
  end else begin
    dat_pre_data[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[50] | in_dat_nan[25])) == 1'b1) begin
    dat_pre_data[407:400] <= dat_pre_data_w[407:400];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[50] | in_dat_nan[25])) == 1'b0) begin
  end else begin
    dat_pre_data[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[51] | in_dat_nan[25])) == 1'b1) begin
    dat_pre_data[415:408] <= dat_pre_data_w[415:408];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[51] | in_dat_nan[25])) == 1'b0) begin
  end else begin
    dat_pre_data[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[52] | in_dat_nan[26])) == 1'b1) begin
    dat_pre_data[423:416] <= dat_pre_data_w[423:416];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[52] | in_dat_nan[26])) == 1'b0) begin
  end else begin
    dat_pre_data[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[53] | in_dat_nan[26])) == 1'b1) begin
    dat_pre_data[431:424] <= dat_pre_data_w[431:424];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[53] | in_dat_nan[26])) == 1'b0) begin
  end else begin
    dat_pre_data[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[54] | in_dat_nan[27])) == 1'b1) begin
    dat_pre_data[439:432] <= dat_pre_data_w[439:432];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[54] | in_dat_nan[27])) == 1'b0) begin
  end else begin
    dat_pre_data[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[55] | in_dat_nan[27])) == 1'b1) begin
    dat_pre_data[447:440] <= dat_pre_data_w[447:440];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[55] | in_dat_nan[27])) == 1'b0) begin
  end else begin
    dat_pre_data[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[56] | in_dat_nan[28])) == 1'b1) begin
    dat_pre_data[455:448] <= dat_pre_data_w[455:448];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[56] | in_dat_nan[28])) == 1'b0) begin
  end else begin
    dat_pre_data[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[57] | in_dat_nan[28])) == 1'b1) begin
    dat_pre_data[463:456] <= dat_pre_data_w[463:456];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[57] | in_dat_nan[28])) == 1'b0) begin
  end else begin
    dat_pre_data[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[58] | in_dat_nan[29])) == 1'b1) begin
    dat_pre_data[471:464] <= dat_pre_data_w[471:464];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[58] | in_dat_nan[29])) == 1'b0) begin
  end else begin
    dat_pre_data[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[59] | in_dat_nan[29])) == 1'b1) begin
    dat_pre_data[479:472] <= dat_pre_data_w[479:472];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[59] | in_dat_nan[29])) == 1'b0) begin
  end else begin
    dat_pre_data[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[60] | in_dat_nan[30])) == 1'b1) begin
    dat_pre_data[487:480] <= dat_pre_data_w[487:480];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[60] | in_dat_nan[30])) == 1'b0) begin
  end else begin
    dat_pre_data[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[61] | in_dat_nan[30])) == 1'b1) begin
    dat_pre_data[495:488] <= dat_pre_data_w[495:488];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[61] | in_dat_nan[30])) == 1'b0) begin
  end else begin
    dat_pre_data[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[62] | in_dat_nan[31])) == 1'b1) begin
    dat_pre_data[503:496] <= dat_pre_data_w[503:496];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[62] | in_dat_nan[31])) == 1'b0) begin
  end else begin
    dat_pre_data[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[63] | in_dat_nan[31])) == 1'b1) begin
    dat_pre_data[511:504] <= dat_pre_data_w[511:504];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[63] | in_dat_nan[31])) == 1'b0) begin
  end else begin
    dat_pre_data[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[64] | in_dat_nan[32])) == 1'b1) begin
    dat_pre_data[519:512] <= dat_pre_data_w[519:512];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[64] | in_dat_nan[32])) == 1'b0) begin
  end else begin
    dat_pre_data[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[65] | in_dat_nan[32])) == 1'b1) begin
    dat_pre_data[527:520] <= dat_pre_data_w[527:520];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[65] | in_dat_nan[32])) == 1'b0) begin
  end else begin
    dat_pre_data[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[66] | in_dat_nan[33])) == 1'b1) begin
    dat_pre_data[535:528] <= dat_pre_data_w[535:528];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[66] | in_dat_nan[33])) == 1'b0) begin
  end else begin
    dat_pre_data[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[67] | in_dat_nan[33])) == 1'b1) begin
    dat_pre_data[543:536] <= dat_pre_data_w[543:536];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[67] | in_dat_nan[33])) == 1'b0) begin
  end else begin
    dat_pre_data[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[68] | in_dat_nan[34])) == 1'b1) begin
    dat_pre_data[551:544] <= dat_pre_data_w[551:544];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[68] | in_dat_nan[34])) == 1'b0) begin
  end else begin
    dat_pre_data[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[69] | in_dat_nan[34])) == 1'b1) begin
    dat_pre_data[559:552] <= dat_pre_data_w[559:552];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[69] | in_dat_nan[34])) == 1'b0) begin
  end else begin
    dat_pre_data[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[70] | in_dat_nan[35])) == 1'b1) begin
    dat_pre_data[567:560] <= dat_pre_data_w[567:560];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[70] | in_dat_nan[35])) == 1'b0) begin
  end else begin
    dat_pre_data[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[71] | in_dat_nan[35])) == 1'b1) begin
    dat_pre_data[575:568] <= dat_pre_data_w[575:568];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[71] | in_dat_nan[35])) == 1'b0) begin
  end else begin
    dat_pre_data[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[72] | in_dat_nan[36])) == 1'b1) begin
    dat_pre_data[583:576] <= dat_pre_data_w[583:576];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[72] | in_dat_nan[36])) == 1'b0) begin
  end else begin
    dat_pre_data[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[73] | in_dat_nan[36])) == 1'b1) begin
    dat_pre_data[591:584] <= dat_pre_data_w[591:584];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[73] | in_dat_nan[36])) == 1'b0) begin
  end else begin
    dat_pre_data[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[74] | in_dat_nan[37])) == 1'b1) begin
    dat_pre_data[599:592] <= dat_pre_data_w[599:592];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[74] | in_dat_nan[37])) == 1'b0) begin
  end else begin
    dat_pre_data[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[75] | in_dat_nan[37])) == 1'b1) begin
    dat_pre_data[607:600] <= dat_pre_data_w[607:600];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[75] | in_dat_nan[37])) == 1'b0) begin
  end else begin
    dat_pre_data[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[76] | in_dat_nan[38])) == 1'b1) begin
    dat_pre_data[615:608] <= dat_pre_data_w[615:608];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[76] | in_dat_nan[38])) == 1'b0) begin
  end else begin
    dat_pre_data[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[77] | in_dat_nan[38])) == 1'b1) begin
    dat_pre_data[623:616] <= dat_pre_data_w[623:616];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[77] | in_dat_nan[38])) == 1'b0) begin
  end else begin
    dat_pre_data[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[78] | in_dat_nan[39])) == 1'b1) begin
    dat_pre_data[631:624] <= dat_pre_data_w[631:624];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[78] | in_dat_nan[39])) == 1'b0) begin
  end else begin
    dat_pre_data[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[79] | in_dat_nan[39])) == 1'b1) begin
    dat_pre_data[639:632] <= dat_pre_data_w[639:632];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[79] | in_dat_nan[39])) == 1'b0) begin
  end else begin
    dat_pre_data[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[80] | in_dat_nan[40])) == 1'b1) begin
    dat_pre_data[647:640] <= dat_pre_data_w[647:640];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[80] | in_dat_nan[40])) == 1'b0) begin
  end else begin
    dat_pre_data[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[81] | in_dat_nan[40])) == 1'b1) begin
    dat_pre_data[655:648] <= dat_pre_data_w[655:648];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[81] | in_dat_nan[40])) == 1'b0) begin
  end else begin
    dat_pre_data[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[82] | in_dat_nan[41])) == 1'b1) begin
    dat_pre_data[663:656] <= dat_pre_data_w[663:656];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[82] | in_dat_nan[41])) == 1'b0) begin
  end else begin
    dat_pre_data[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[83] | in_dat_nan[41])) == 1'b1) begin
    dat_pre_data[671:664] <= dat_pre_data_w[671:664];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[83] | in_dat_nan[41])) == 1'b0) begin
  end else begin
    dat_pre_data[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[84] | in_dat_nan[42])) == 1'b1) begin
    dat_pre_data[679:672] <= dat_pre_data_w[679:672];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[84] | in_dat_nan[42])) == 1'b0) begin
  end else begin
    dat_pre_data[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[85] | in_dat_nan[42])) == 1'b1) begin
    dat_pre_data[687:680] <= dat_pre_data_w[687:680];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[85] | in_dat_nan[42])) == 1'b0) begin
  end else begin
    dat_pre_data[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[86] | in_dat_nan[43])) == 1'b1) begin
    dat_pre_data[695:688] <= dat_pre_data_w[695:688];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[86] | in_dat_nan[43])) == 1'b0) begin
  end else begin
    dat_pre_data[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[87] | in_dat_nan[43])) == 1'b1) begin
    dat_pre_data[703:696] <= dat_pre_data_w[703:696];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[87] | in_dat_nan[43])) == 1'b0) begin
  end else begin
    dat_pre_data[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[88] | in_dat_nan[44])) == 1'b1) begin
    dat_pre_data[711:704] <= dat_pre_data_w[711:704];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[88] | in_dat_nan[44])) == 1'b0) begin
  end else begin
    dat_pre_data[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[89] | in_dat_nan[44])) == 1'b1) begin
    dat_pre_data[719:712] <= dat_pre_data_w[719:712];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[89] | in_dat_nan[44])) == 1'b0) begin
  end else begin
    dat_pre_data[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[90] | in_dat_nan[45])) == 1'b1) begin
    dat_pre_data[727:720] <= dat_pre_data_w[727:720];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[90] | in_dat_nan[45])) == 1'b0) begin
  end else begin
    dat_pre_data[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[91] | in_dat_nan[45])) == 1'b1) begin
    dat_pre_data[735:728] <= dat_pre_data_w[735:728];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[91] | in_dat_nan[45])) == 1'b0) begin
  end else begin
    dat_pre_data[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[92] | in_dat_nan[46])) == 1'b1) begin
    dat_pre_data[743:736] <= dat_pre_data_w[743:736];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[92] | in_dat_nan[46])) == 1'b0) begin
  end else begin
    dat_pre_data[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[93] | in_dat_nan[46])) == 1'b1) begin
    dat_pre_data[751:744] <= dat_pre_data_w[751:744];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[93] | in_dat_nan[46])) == 1'b0) begin
  end else begin
    dat_pre_data[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[94] | in_dat_nan[47])) == 1'b1) begin
    dat_pre_data[759:752] <= dat_pre_data_w[759:752];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[94] | in_dat_nan[47])) == 1'b0) begin
  end else begin
    dat_pre_data[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[95] | in_dat_nan[47])) == 1'b1) begin
    dat_pre_data[767:760] <= dat_pre_data_w[767:760];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[95] | in_dat_nan[47])) == 1'b0) begin
  end else begin
    dat_pre_data[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[96] | in_dat_nan[48])) == 1'b1) begin
    dat_pre_data[775:768] <= dat_pre_data_w[775:768];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[96] | in_dat_nan[48])) == 1'b0) begin
  end else begin
    dat_pre_data[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[97] | in_dat_nan[48])) == 1'b1) begin
    dat_pre_data[783:776] <= dat_pre_data_w[783:776];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[97] | in_dat_nan[48])) == 1'b0) begin
  end else begin
    dat_pre_data[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[98] | in_dat_nan[49])) == 1'b1) begin
    dat_pre_data[791:784] <= dat_pre_data_w[791:784];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[98] | in_dat_nan[49])) == 1'b0) begin
  end else begin
    dat_pre_data[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[99] | in_dat_nan[49])) == 1'b1) begin
    dat_pre_data[799:792] <= dat_pre_data_w[799:792];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[99] | in_dat_nan[49])) == 1'b0) begin
  end else begin
    dat_pre_data[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[100] | in_dat_nan[50])) == 1'b1) begin
    dat_pre_data[807:800] <= dat_pre_data_w[807:800];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[100] | in_dat_nan[50])) == 1'b0) begin
  end else begin
    dat_pre_data[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[101] | in_dat_nan[50])) == 1'b1) begin
    dat_pre_data[815:808] <= dat_pre_data_w[815:808];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[101] | in_dat_nan[50])) == 1'b0) begin
  end else begin
    dat_pre_data[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[102] | in_dat_nan[51])) == 1'b1) begin
    dat_pre_data[823:816] <= dat_pre_data_w[823:816];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[102] | in_dat_nan[51])) == 1'b0) begin
  end else begin
    dat_pre_data[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[103] | in_dat_nan[51])) == 1'b1) begin
    dat_pre_data[831:824] <= dat_pre_data_w[831:824];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[103] | in_dat_nan[51])) == 1'b0) begin
  end else begin
    dat_pre_data[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[104] | in_dat_nan[52])) == 1'b1) begin
    dat_pre_data[839:832] <= dat_pre_data_w[839:832];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[104] | in_dat_nan[52])) == 1'b0) begin
  end else begin
    dat_pre_data[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[105] | in_dat_nan[52])) == 1'b1) begin
    dat_pre_data[847:840] <= dat_pre_data_w[847:840];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[105] | in_dat_nan[52])) == 1'b0) begin
  end else begin
    dat_pre_data[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[106] | in_dat_nan[53])) == 1'b1) begin
    dat_pre_data[855:848] <= dat_pre_data_w[855:848];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[106] | in_dat_nan[53])) == 1'b0) begin
  end else begin
    dat_pre_data[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[107] | in_dat_nan[53])) == 1'b1) begin
    dat_pre_data[863:856] <= dat_pre_data_w[863:856];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[107] | in_dat_nan[53])) == 1'b0) begin
  end else begin
    dat_pre_data[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[108] | in_dat_nan[54])) == 1'b1) begin
    dat_pre_data[871:864] <= dat_pre_data_w[871:864];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[108] | in_dat_nan[54])) == 1'b0) begin
  end else begin
    dat_pre_data[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[109] | in_dat_nan[54])) == 1'b1) begin
    dat_pre_data[879:872] <= dat_pre_data_w[879:872];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[109] | in_dat_nan[54])) == 1'b0) begin
  end else begin
    dat_pre_data[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[110] | in_dat_nan[55])) == 1'b1) begin
    dat_pre_data[887:880] <= dat_pre_data_w[887:880];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[110] | in_dat_nan[55])) == 1'b0) begin
  end else begin
    dat_pre_data[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[111] | in_dat_nan[55])) == 1'b1) begin
    dat_pre_data[895:888] <= dat_pre_data_w[895:888];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[111] | in_dat_nan[55])) == 1'b0) begin
  end else begin
    dat_pre_data[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[112] | in_dat_nan[56])) == 1'b1) begin
    dat_pre_data[903:896] <= dat_pre_data_w[903:896];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[112] | in_dat_nan[56])) == 1'b0) begin
  end else begin
    dat_pre_data[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[113] | in_dat_nan[56])) == 1'b1) begin
    dat_pre_data[911:904] <= dat_pre_data_w[911:904];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[113] | in_dat_nan[56])) == 1'b0) begin
  end else begin
    dat_pre_data[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[114] | in_dat_nan[57])) == 1'b1) begin
    dat_pre_data[919:912] <= dat_pre_data_w[919:912];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[114] | in_dat_nan[57])) == 1'b0) begin
  end else begin
    dat_pre_data[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[115] | in_dat_nan[57])) == 1'b1) begin
    dat_pre_data[927:920] <= dat_pre_data_w[927:920];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[115] | in_dat_nan[57])) == 1'b0) begin
  end else begin
    dat_pre_data[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[116] | in_dat_nan[58])) == 1'b1) begin
    dat_pre_data[935:928] <= dat_pre_data_w[935:928];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[116] | in_dat_nan[58])) == 1'b0) begin
  end else begin
    dat_pre_data[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[117] | in_dat_nan[58])) == 1'b1) begin
    dat_pre_data[943:936] <= dat_pre_data_w[943:936];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[117] | in_dat_nan[58])) == 1'b0) begin
  end else begin
    dat_pre_data[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[118] | in_dat_nan[59])) == 1'b1) begin
    dat_pre_data[951:944] <= dat_pre_data_w[951:944];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[118] | in_dat_nan[59])) == 1'b0) begin
  end else begin
    dat_pre_data[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[119] | in_dat_nan[59])) == 1'b1) begin
    dat_pre_data[959:952] <= dat_pre_data_w[959:952];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[119] | in_dat_nan[59])) == 1'b0) begin
  end else begin
    dat_pre_data[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[120] | in_dat_nan[60])) == 1'b1) begin
    dat_pre_data[967:960] <= dat_pre_data_w[967:960];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[120] | in_dat_nan[60])) == 1'b0) begin
  end else begin
    dat_pre_data[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[121] | in_dat_nan[60])) == 1'b1) begin
    dat_pre_data[975:968] <= dat_pre_data_w[975:968];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[121] | in_dat_nan[60])) == 1'b0) begin
  end else begin
    dat_pre_data[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[122] | in_dat_nan[61])) == 1'b1) begin
    dat_pre_data[983:976] <= dat_pre_data_w[983:976];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[122] | in_dat_nan[61])) == 1'b0) begin
  end else begin
    dat_pre_data[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[123] | in_dat_nan[61])) == 1'b1) begin
    dat_pre_data[991:984] <= dat_pre_data_w[991:984];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[123] | in_dat_nan[61])) == 1'b0) begin
  end else begin
    dat_pre_data[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[124] | in_dat_nan[62])) == 1'b1) begin
    dat_pre_data[999:992] <= dat_pre_data_w[999:992];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[124] | in_dat_nan[62])) == 1'b0) begin
  end else begin
    dat_pre_data[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[125] | in_dat_nan[62])) == 1'b1) begin
    dat_pre_data[1007:1000] <= dat_pre_data_w[1007:1000];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[125] | in_dat_nan[62])) == 1'b0) begin
  end else begin
    dat_pre_data[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[126] | in_dat_nan[63])) == 1'b1) begin
    dat_pre_data[1015:1008] <= dat_pre_data_w[1015:1008];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[126] | in_dat_nan[63])) == 1'b0) begin
  end else begin
    dat_pre_data[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & (dat_pre_nz_w[127] | in_dat_nan[63])) == 1'b1) begin
    dat_pre_data[1023:1016] <= dat_pre_data_w[1023:1016];
  // VCS coverage off
  end else if ((in_dat_pvld & (dat_pre_nz_w[127] | in_dat_nan[63])) == 1'b0) begin
  end else begin
    dat_pre_data[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_pre_stripe_st <= {16{1'b0}};
  end else begin
  dat_pre_stripe_st <= {16{in_dat_stripe_st & in_dat_pvld}};
  end
end
always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_pre_stripe_end <= {9{1'b0}};
  end else begin
  dat_pre_stripe_end <= {9{in_dat_stripe_end & in_dat_pvld}};
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[82]) == 1'b1) begin
    dat_pre_mask0 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[82]) == 1'b0) begin
  end else begin
    dat_pre_mask0 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[82]) == 1'b1) begin
    dat_pre_exp_reg0 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[82]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg0 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[83]) == 1'b1) begin
    dat_pre_mask1 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[83]) == 1'b0) begin
  end else begin
    dat_pre_mask1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[83]) == 1'b1) begin
    dat_pre_exp_reg1 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[83]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[84]) == 1'b1) begin
    dat_pre_mask2 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[84]) == 1'b0) begin
  end else begin
    dat_pre_mask2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[84]) == 1'b1) begin
    dat_pre_exp_reg2 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[84]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[85]) == 1'b1) begin
    dat_pre_mask3 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[85]) == 1'b0) begin
  end else begin
    dat_pre_mask3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[85]) == 1'b1) begin
    dat_pre_exp_reg3 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[85]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[86]) == 1'b1) begin
    dat_pre_mask4 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[86]) == 1'b0) begin
  end else begin
    dat_pre_mask4 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[86]) == 1'b1) begin
    dat_pre_exp_reg4 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[86]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg4 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[87]) == 1'b1) begin
    dat_pre_mask5 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[87]) == 1'b0) begin
  end else begin
    dat_pre_mask5 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[87]) == 1'b1) begin
    dat_pre_exp_reg5 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[87]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg5 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[88]) == 1'b1) begin
    dat_pre_mask6 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[88]) == 1'b0) begin
  end else begin
    dat_pre_mask6 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[88]) == 1'b1) begin
    dat_pre_exp_reg6 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[88]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg6 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end


always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[89]) == 1'b1) begin
    dat_pre_mask7 <= dat_pre_mask_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[89]) == 1'b0) begin
  end else begin
    dat_pre_mask7 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((in_dat_pvld & cfg_is_fp16_d1[89]) == 1'b1) begin
    dat_pre_exp_reg7 <= dat_pre_exp_w;
  // VCS coverage off
  end else if ((in_dat_pvld & cfg_is_fp16_d1[89]) == 1'b0) begin
  end else begin
    dat_pre_exp_reg7 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end





always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask0
  or dat_pre_exp_reg0
  ) begin
    dat0_pre_pvld       = dat_pre_pvld[0];
    dat0_pre_stripe_st  = dat_pre_stripe_st[0+8];
    dat0_pre_stripe_end = dat_pre_stripe_end[0];
    dat0_pre_mask       = dat_pre_mask0;
    dat0_pre_exp        = dat_pre_exp_reg0;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask1
  or dat_pre_exp_reg1
  ) begin
    dat1_pre_pvld       = dat_pre_pvld[1];
    dat1_pre_stripe_st  = dat_pre_stripe_st[1+8];
    dat1_pre_stripe_end = dat_pre_stripe_end[1];
    dat1_pre_mask       = dat_pre_mask1;
    dat1_pre_exp        = dat_pre_exp_reg1;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask2
  or dat_pre_exp_reg2
  ) begin
    dat2_pre_pvld       = dat_pre_pvld[2];
    dat2_pre_stripe_st  = dat_pre_stripe_st[2+8];
    dat2_pre_stripe_end = dat_pre_stripe_end[2];
    dat2_pre_mask       = dat_pre_mask2;
    dat2_pre_exp        = dat_pre_exp_reg2;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask3
  or dat_pre_exp_reg3
  ) begin
    dat3_pre_pvld       = dat_pre_pvld[3];
    dat3_pre_stripe_st  = dat_pre_stripe_st[3+8];
    dat3_pre_stripe_end = dat_pre_stripe_end[3];
    dat3_pre_mask       = dat_pre_mask3;
    dat3_pre_exp        = dat_pre_exp_reg3;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask4
  or dat_pre_exp_reg4
  ) begin
    dat4_pre_pvld       = dat_pre_pvld[4];
    dat4_pre_stripe_st  = dat_pre_stripe_st[4+8];
    dat4_pre_stripe_end = dat_pre_stripe_end[4];
    dat4_pre_mask       = dat_pre_mask4;
    dat4_pre_exp        = dat_pre_exp_reg4;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask5
  or dat_pre_exp_reg5
  ) begin
    dat5_pre_pvld       = dat_pre_pvld[5];
    dat5_pre_stripe_st  = dat_pre_stripe_st[5+8];
    dat5_pre_stripe_end = dat_pre_stripe_end[5];
    dat5_pre_mask       = dat_pre_mask5;
    dat5_pre_exp        = dat_pre_exp_reg5;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask6
  or dat_pre_exp_reg6
  ) begin
    dat6_pre_pvld       = dat_pre_pvld[6];
    dat6_pre_stripe_st  = dat_pre_stripe_st[6+8];
    dat6_pre_stripe_end = dat_pre_stripe_end[6];
    dat6_pre_mask       = dat_pre_mask6;
    dat6_pre_exp        = dat_pre_exp_reg6;
end


always @(
  dat_pre_pvld
  or dat_pre_stripe_st
  or dat_pre_stripe_end
  or dat_pre_mask7
  or dat_pre_exp_reg7
  ) begin
    dat7_pre_pvld       = dat_pre_pvld[7];
    dat7_pre_stripe_st  = dat_pre_stripe_st[7+8];
    dat7_pre_stripe_end = dat_pre_stripe_end[7];
    dat7_pre_mask       = dat_pre_mask7;
    dat7_pre_exp        = dat_pre_exp_reg7;
end





//==========================================================
// Data active register         
//==========================================================

always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg0 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg0 <= {104{dat_pre_pvld[8]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8]) == 1'b1) begin
    dat_actv_nz_reg0 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[8]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg0 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & cfg_is_fp16_d1[90]) == 1'b1) begin
    dat_actv_nan_reg0 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & cfg_is_fp16_d1[90]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg0 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg0[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg0[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg0[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg0[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg0[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg0[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg0[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg0[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg0[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg0[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg0[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg0[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg0[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg0[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg0[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg0[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg0[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg0[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg0[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg0[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg0[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg0[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg0[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg0[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg0[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg0[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg0[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg0[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg0[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg0[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg0[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg0[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg0[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg0[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg0[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg0[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg0[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg0[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg0[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg0[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg0[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg0[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg0[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg0[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg0[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg0[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg0[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg0[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg0[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg0[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg0[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg0[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg0[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg0[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg0[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg0[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg0[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg0[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg0[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg0[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg0[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg0[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg0[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg0[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg0[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg0[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg0[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg0[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg0[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg0[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg0[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg0[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg0[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg0[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg0[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg0[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg0[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg0[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg0[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg0[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg0[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg0[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg0[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg0[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg0[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg0[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg0[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg0[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg0[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg0[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg0[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg0[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg0[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg0[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg0[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg0[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg0[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg0[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg0[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg0[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg0[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg0[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg0[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg0[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg0[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg0[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg0[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg0[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg0[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg0[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg0[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg0[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg0[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg0[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg0[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg0[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg0[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg0[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg0[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg0[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg0[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg0[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg0[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg0[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg0[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg0[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg0[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[8] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg0[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[8] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg0[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg1 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg1 <= {104{dat_pre_pvld[9]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9]) == 1'b1) begin
    dat_actv_nz_reg1 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[9]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & cfg_is_fp16_d1[91]) == 1'b1) begin
    dat_actv_nan_reg1 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & cfg_is_fp16_d1[91]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg1 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg1[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg1[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg1[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg1[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg1[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg1[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg1[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg1[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg1[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg1[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg1[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg1[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg1[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg1[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg1[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg1[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg1[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg1[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg1[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg1[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg1[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg1[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg1[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg1[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg1[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg1[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg1[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg1[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg1[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg1[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg1[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg1[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg1[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg1[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg1[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg1[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg1[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg1[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg1[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg1[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg1[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg1[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg1[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg1[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg1[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg1[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg1[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg1[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg1[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg1[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg1[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg1[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg1[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg1[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg1[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg1[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg1[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg1[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg1[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg1[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg1[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg1[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg1[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg1[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg1[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg1[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg1[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg1[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg1[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg1[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg1[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg1[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg1[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg1[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg1[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg1[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg1[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg1[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg1[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg1[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg1[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg1[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg1[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg1[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg1[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg1[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg1[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg1[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg1[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg1[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg1[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg1[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg1[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg1[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg1[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg1[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg1[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg1[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg1[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg1[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg1[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg1[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg1[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg1[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg1[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg1[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg1[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg1[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg1[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg1[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg1[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg1[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg1[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg1[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg1[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg1[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg1[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg1[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg1[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg1[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg1[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg1[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg1[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg1[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg1[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg1[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg1[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[9] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg1[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[9] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg1[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg2 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg2 <= {104{dat_pre_pvld[10]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10]) == 1'b1) begin
    dat_actv_nz_reg2 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[10]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & cfg_is_fp16_d1[92]) == 1'b1) begin
    dat_actv_nan_reg2 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & cfg_is_fp16_d1[92]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg2 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg2[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg2[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg2[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg2[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg2[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg2[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg2[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg2[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg2[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg2[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg2[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg2[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg2[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg2[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg2[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg2[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg2[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg2[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg2[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg2[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg2[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg2[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg2[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg2[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg2[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg2[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg2[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg2[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg2[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg2[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg2[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg2[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg2[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg2[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg2[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg2[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg2[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg2[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg2[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg2[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg2[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg2[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg2[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg2[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg2[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg2[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg2[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg2[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg2[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg2[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg2[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg2[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg2[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg2[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg2[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg2[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg2[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg2[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg2[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg2[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg2[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg2[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg2[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg2[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg2[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg2[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg2[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg2[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg2[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg2[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg2[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg2[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg2[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg2[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg2[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg2[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg2[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg2[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg2[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg2[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg2[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg2[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg2[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg2[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg2[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg2[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg2[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg2[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg2[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg2[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg2[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg2[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg2[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg2[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg2[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg2[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg2[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg2[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg2[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg2[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg2[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg2[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg2[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg2[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg2[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg2[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg2[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg2[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg2[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg2[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg2[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg2[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg2[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg2[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg2[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg2[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg2[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg2[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg2[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg2[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg2[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg2[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg2[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg2[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg2[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg2[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg2[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[10] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg2[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[10] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg2[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg3 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg3 <= {104{dat_pre_pvld[11]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11]) == 1'b1) begin
    dat_actv_nz_reg3 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[11]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & cfg_is_fp16_d1[93]) == 1'b1) begin
    dat_actv_nan_reg3 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & cfg_is_fp16_d1[93]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg3 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg3[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg3[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg3[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg3[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg3[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg3[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg3[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg3[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg3[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg3[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg3[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg3[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg3[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg3[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg3[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg3[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg3[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg3[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg3[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg3[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg3[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg3[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg3[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg3[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg3[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg3[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg3[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg3[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg3[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg3[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg3[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg3[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg3[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg3[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg3[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg3[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg3[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg3[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg3[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg3[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg3[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg3[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg3[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg3[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg3[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg3[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg3[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg3[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg3[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg3[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg3[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg3[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg3[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg3[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg3[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg3[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg3[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg3[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg3[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg3[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg3[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg3[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg3[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg3[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg3[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg3[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg3[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg3[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg3[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg3[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg3[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg3[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg3[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg3[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg3[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg3[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg3[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg3[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg3[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg3[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg3[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg3[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg3[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg3[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg3[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg3[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg3[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg3[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg3[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg3[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg3[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg3[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg3[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg3[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg3[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg3[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg3[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg3[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg3[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg3[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg3[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg3[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg3[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg3[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg3[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg3[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg3[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg3[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg3[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg3[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg3[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg3[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg3[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg3[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg3[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg3[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg3[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg3[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg3[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg3[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg3[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg3[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg3[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg3[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg3[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg3[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg3[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[11] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg3[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[11] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg3[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg4 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg4 <= {104{dat_pre_pvld[12]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12]) == 1'b1) begin
    dat_actv_nz_reg4 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[12]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg4 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & cfg_is_fp16_d1[94]) == 1'b1) begin
    dat_actv_nan_reg4 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & cfg_is_fp16_d1[94]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg4 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg4[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg4[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg4[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg4[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg4[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg4[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg4[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg4[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg4[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg4[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg4[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg4[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg4[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg4[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg4[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg4[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg4[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg4[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg4[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg4[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg4[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg4[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg4[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg4[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg4[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg4[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg4[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg4[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg4[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg4[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg4[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg4[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg4[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg4[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg4[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg4[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg4[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg4[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg4[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg4[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg4[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg4[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg4[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg4[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg4[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg4[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg4[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg4[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg4[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg4[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg4[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg4[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg4[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg4[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg4[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg4[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg4[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg4[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg4[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg4[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg4[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg4[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg4[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg4[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg4[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg4[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg4[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg4[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg4[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg4[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg4[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg4[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg4[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg4[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg4[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg4[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg4[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg4[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg4[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg4[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg4[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg4[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg4[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg4[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg4[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg4[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg4[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg4[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg4[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg4[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg4[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg4[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg4[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg4[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg4[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg4[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg4[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg4[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg4[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg4[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg4[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg4[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg4[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg4[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg4[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg4[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg4[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg4[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg4[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg4[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg4[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg4[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg4[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg4[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg4[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg4[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg4[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg4[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg4[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg4[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg4[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg4[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg4[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg4[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg4[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg4[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg4[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[12] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg4[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[12] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg4[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg5 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg5 <= {104{dat_pre_pvld[13]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13]) == 1'b1) begin
    dat_actv_nz_reg5 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[13]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg5 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & cfg_is_fp16_d1[95]) == 1'b1) begin
    dat_actv_nan_reg5 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & cfg_is_fp16_d1[95]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg5 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg5[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg5[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg5[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg5[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg5[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg5[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg5[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg5[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg5[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg5[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg5[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg5[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg5[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg5[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg5[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg5[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg5[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg5[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg5[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg5[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg5[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg5[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg5[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg5[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg5[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg5[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg5[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg5[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg5[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg5[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg5[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg5[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg5[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg5[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg5[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg5[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg5[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg5[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg5[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg5[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg5[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg5[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg5[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg5[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg5[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg5[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg5[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg5[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg5[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg5[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg5[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg5[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg5[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg5[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg5[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg5[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg5[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg5[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg5[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg5[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg5[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg5[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg5[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg5[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg5[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg5[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg5[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg5[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg5[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg5[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg5[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg5[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg5[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg5[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg5[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg5[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg5[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg5[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg5[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg5[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg5[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg5[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg5[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg5[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg5[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg5[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg5[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg5[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg5[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg5[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg5[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg5[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg5[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg5[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg5[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg5[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg5[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg5[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg5[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg5[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg5[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg5[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg5[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg5[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg5[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg5[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg5[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg5[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg5[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg5[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg5[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg5[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg5[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg5[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg5[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg5[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg5[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg5[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg5[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg5[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg5[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg5[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg5[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg5[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg5[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg5[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg5[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[13] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg5[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[13] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg5[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg6 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg6 <= {104{dat_pre_pvld[14]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14]) == 1'b1) begin
    dat_actv_nz_reg6 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[14]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg6 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & cfg_is_fp16_d1[96]) == 1'b1) begin
    dat_actv_nan_reg6 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & cfg_is_fp16_d1[96]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg6 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg6[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg6[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg6[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg6[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg6[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg6[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg6[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg6[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg6[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg6[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg6[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg6[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg6[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg6[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg6[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg6[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg6[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg6[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg6[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg6[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg6[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg6[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg6[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg6[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg6[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg6[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg6[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg6[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg6[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg6[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg6[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg6[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg6[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg6[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg6[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg6[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg6[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg6[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg6[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg6[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg6[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg6[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg6[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg6[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg6[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg6[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg6[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg6[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg6[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg6[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg6[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg6[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg6[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg6[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg6[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg6[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg6[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg6[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg6[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg6[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg6[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg6[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg6[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg6[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg6[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg6[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg6[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg6[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg6[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg6[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg6[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg6[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg6[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg6[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg6[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg6[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg6[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg6[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg6[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg6[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg6[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg6[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg6[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg6[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg6[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg6[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg6[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg6[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg6[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg6[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg6[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg6[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg6[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg6[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg6[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg6[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg6[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg6[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg6[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg6[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg6[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg6[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg6[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg6[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg6[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg6[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg6[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg6[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg6[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg6[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg6[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg6[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg6[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg6[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg6[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg6[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg6[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg6[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg6[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg6[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg6[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg6[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg6[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg6[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg6[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg6[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg6[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[14] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg6[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[14] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg6[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end




always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
  if (!nvdla_core_rstn) begin
    dat_actv_pvld_reg7 <= {104{1'b0}};
  end else begin
  dat_actv_pvld_reg7 <= {104{dat_pre_pvld[15]}};
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15]) == 1'b1) begin
    dat_actv_nz_reg7 <= dat_pre_nz;
  // VCS coverage off
  end else if ((dat_pre_pvld[15]) == 1'b0) begin
  end else begin
    dat_actv_nz_reg7 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & cfg_is_fp16_d1[97]) == 1'b1) begin
    dat_actv_nan_reg7 <= dat_pre_nan;
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & cfg_is_fp16_d1[97]) == 1'b0) begin
  end else begin
    dat_actv_nan_reg7 <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end

always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg7[7:0] <= dat_pre_data[7:0];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[0] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[7:0] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b1) begin
    dat_actv_data_reg7[15:8] <= dat_pre_data[15:8];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[1] | dat_pre_nan[0])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[15:8] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg7[23:16] <= dat_pre_data[23:16];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[2] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[23:16] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b1) begin
    dat_actv_data_reg7[31:24] <= dat_pre_data[31:24];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[3] | dat_pre_nan[1])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[31:24] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg7[39:32] <= dat_pre_data[39:32];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[4] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[39:32] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b1) begin
    dat_actv_data_reg7[47:40] <= dat_pre_data[47:40];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[5] | dat_pre_nan[2])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[47:40] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg7[55:48] <= dat_pre_data[55:48];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[6] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[55:48] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b1) begin
    dat_actv_data_reg7[63:56] <= dat_pre_data[63:56];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[7] | dat_pre_nan[3])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[63:56] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg7[71:64] <= dat_pre_data[71:64];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[8] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[71:64] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b1) begin
    dat_actv_data_reg7[79:72] <= dat_pre_data[79:72];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[9] | dat_pre_nan[4])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[79:72] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg7[87:80] <= dat_pre_data[87:80];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[10] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[87:80] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b1) begin
    dat_actv_data_reg7[95:88] <= dat_pre_data[95:88];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[11] | dat_pre_nan[5])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[95:88] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg7[103:96] <= dat_pre_data[103:96];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[12] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[103:96] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b1) begin
    dat_actv_data_reg7[111:104] <= dat_pre_data[111:104];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[13] | dat_pre_nan[6])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[111:104] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg7[119:112] <= dat_pre_data[119:112];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[14] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[119:112] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b1) begin
    dat_actv_data_reg7[127:120] <= dat_pre_data[127:120];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[15] | dat_pre_nan[7])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[127:120] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg7[135:128] <= dat_pre_data[135:128];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[16] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[135:128] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b1) begin
    dat_actv_data_reg7[143:136] <= dat_pre_data[143:136];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[17] | dat_pre_nan[8])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[143:136] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg7[151:144] <= dat_pre_data[151:144];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[18] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[151:144] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b1) begin
    dat_actv_data_reg7[159:152] <= dat_pre_data[159:152];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[19] | dat_pre_nan[9])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[159:152] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg7[167:160] <= dat_pre_data[167:160];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[20] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[167:160] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b1) begin
    dat_actv_data_reg7[175:168] <= dat_pre_data[175:168];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[21] | dat_pre_nan[10])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[175:168] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg7[183:176] <= dat_pre_data[183:176];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[22] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[183:176] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b1) begin
    dat_actv_data_reg7[191:184] <= dat_pre_data[191:184];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[23] | dat_pre_nan[11])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[191:184] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg7[199:192] <= dat_pre_data[199:192];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[24] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[199:192] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b1) begin
    dat_actv_data_reg7[207:200] <= dat_pre_data[207:200];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[25] | dat_pre_nan[12])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[207:200] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg7[215:208] <= dat_pre_data[215:208];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[26] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[215:208] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b1) begin
    dat_actv_data_reg7[223:216] <= dat_pre_data[223:216];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[27] | dat_pre_nan[13])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[223:216] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg7[231:224] <= dat_pre_data[231:224];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[28] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[231:224] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b1) begin
    dat_actv_data_reg7[239:232] <= dat_pre_data[239:232];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[29] | dat_pre_nan[14])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[239:232] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg7[247:240] <= dat_pre_data[247:240];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[30] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[247:240] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b1) begin
    dat_actv_data_reg7[255:248] <= dat_pre_data[255:248];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[31] | dat_pre_nan[15])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[255:248] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg7[263:256] <= dat_pre_data[263:256];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[32] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[263:256] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b1) begin
    dat_actv_data_reg7[271:264] <= dat_pre_data[271:264];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[33] | dat_pre_nan[16])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[271:264] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg7[279:272] <= dat_pre_data[279:272];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[34] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[279:272] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b1) begin
    dat_actv_data_reg7[287:280] <= dat_pre_data[287:280];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[35] | dat_pre_nan[17])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[287:280] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg7[295:288] <= dat_pre_data[295:288];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[36] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[295:288] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b1) begin
    dat_actv_data_reg7[303:296] <= dat_pre_data[303:296];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[37] | dat_pre_nan[18])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[303:296] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg7[311:304] <= dat_pre_data[311:304];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[38] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[311:304] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b1) begin
    dat_actv_data_reg7[319:312] <= dat_pre_data[319:312];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[39] | dat_pre_nan[19])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[319:312] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg7[327:320] <= dat_pre_data[327:320];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[40] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[327:320] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b1) begin
    dat_actv_data_reg7[335:328] <= dat_pre_data[335:328];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[41] | dat_pre_nan[20])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[335:328] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg7[343:336] <= dat_pre_data[343:336];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[42] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[343:336] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b1) begin
    dat_actv_data_reg7[351:344] <= dat_pre_data[351:344];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[43] | dat_pre_nan[21])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[351:344] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg7[359:352] <= dat_pre_data[359:352];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[44] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[359:352] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b1) begin
    dat_actv_data_reg7[367:360] <= dat_pre_data[367:360];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[45] | dat_pre_nan[22])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[367:360] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg7[375:368] <= dat_pre_data[375:368];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[46] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[375:368] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b1) begin
    dat_actv_data_reg7[383:376] <= dat_pre_data[383:376];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[47] | dat_pre_nan[23])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[383:376] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg7[391:384] <= dat_pre_data[391:384];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[48] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[391:384] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b1) begin
    dat_actv_data_reg7[399:392] <= dat_pre_data[399:392];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[49] | dat_pre_nan[24])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[399:392] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg7[407:400] <= dat_pre_data[407:400];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[50] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[407:400] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b1) begin
    dat_actv_data_reg7[415:408] <= dat_pre_data[415:408];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[51] | dat_pre_nan[25])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[415:408] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg7[423:416] <= dat_pre_data[423:416];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[52] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[423:416] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b1) begin
    dat_actv_data_reg7[431:424] <= dat_pre_data[431:424];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[53] | dat_pre_nan[26])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[431:424] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg7[439:432] <= dat_pre_data[439:432];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[54] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[439:432] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b1) begin
    dat_actv_data_reg7[447:440] <= dat_pre_data[447:440];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[55] | dat_pre_nan[27])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[447:440] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg7[455:448] <= dat_pre_data[455:448];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[56] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[455:448] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b1) begin
    dat_actv_data_reg7[463:456] <= dat_pre_data[463:456];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[57] | dat_pre_nan[28])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[463:456] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg7[471:464] <= dat_pre_data[471:464];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[58] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[471:464] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b1) begin
    dat_actv_data_reg7[479:472] <= dat_pre_data[479:472];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[59] | dat_pre_nan[29])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[479:472] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg7[487:480] <= dat_pre_data[487:480];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[60] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[487:480] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b1) begin
    dat_actv_data_reg7[495:488] <= dat_pre_data[495:488];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[61] | dat_pre_nan[30])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[495:488] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg7[503:496] <= dat_pre_data[503:496];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[62] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[503:496] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b1) begin
    dat_actv_data_reg7[511:504] <= dat_pre_data[511:504];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[63] | dat_pre_nan[31])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[511:504] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg7[519:512] <= dat_pre_data[519:512];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[64] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[519:512] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b1) begin
    dat_actv_data_reg7[527:520] <= dat_pre_data[527:520];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[65] | dat_pre_nan[32])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[527:520] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg7[535:528] <= dat_pre_data[535:528];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[66] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[535:528] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b1) begin
    dat_actv_data_reg7[543:536] <= dat_pre_data[543:536];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[67] | dat_pre_nan[33])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[543:536] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg7[551:544] <= dat_pre_data[551:544];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[68] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[551:544] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b1) begin
    dat_actv_data_reg7[559:552] <= dat_pre_data[559:552];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[69] | dat_pre_nan[34])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[559:552] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg7[567:560] <= dat_pre_data[567:560];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[70] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[567:560] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b1) begin
    dat_actv_data_reg7[575:568] <= dat_pre_data[575:568];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[71] | dat_pre_nan[35])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[575:568] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg7[583:576] <= dat_pre_data[583:576];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[72] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[583:576] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b1) begin
    dat_actv_data_reg7[591:584] <= dat_pre_data[591:584];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[73] | dat_pre_nan[36])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[591:584] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg7[599:592] <= dat_pre_data[599:592];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[74] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[599:592] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b1) begin
    dat_actv_data_reg7[607:600] <= dat_pre_data[607:600];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[75] | dat_pre_nan[37])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[607:600] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg7[615:608] <= dat_pre_data[615:608];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[76] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[615:608] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b1) begin
    dat_actv_data_reg7[623:616] <= dat_pre_data[623:616];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[77] | dat_pre_nan[38])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[623:616] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg7[631:624] <= dat_pre_data[631:624];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[78] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[631:624] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b1) begin
    dat_actv_data_reg7[639:632] <= dat_pre_data[639:632];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[79] | dat_pre_nan[39])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[639:632] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg7[647:640] <= dat_pre_data[647:640];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[80] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[647:640] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b1) begin
    dat_actv_data_reg7[655:648] <= dat_pre_data[655:648];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[81] | dat_pre_nan[40])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[655:648] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg7[663:656] <= dat_pre_data[663:656];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[82] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[663:656] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b1) begin
    dat_actv_data_reg7[671:664] <= dat_pre_data[671:664];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[83] | dat_pre_nan[41])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[671:664] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg7[679:672] <= dat_pre_data[679:672];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[84] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[679:672] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b1) begin
    dat_actv_data_reg7[687:680] <= dat_pre_data[687:680];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[85] | dat_pre_nan[42])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[687:680] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg7[695:688] <= dat_pre_data[695:688];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[86] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[695:688] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b1) begin
    dat_actv_data_reg7[703:696] <= dat_pre_data[703:696];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[87] | dat_pre_nan[43])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[703:696] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg7[711:704] <= dat_pre_data[711:704];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[88] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[711:704] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b1) begin
    dat_actv_data_reg7[719:712] <= dat_pre_data[719:712];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[89] | dat_pre_nan[44])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[719:712] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg7[727:720] <= dat_pre_data[727:720];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[90] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[727:720] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b1) begin
    dat_actv_data_reg7[735:728] <= dat_pre_data[735:728];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[91] | dat_pre_nan[45])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[735:728] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg7[743:736] <= dat_pre_data[743:736];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[92] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[743:736] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b1) begin
    dat_actv_data_reg7[751:744] <= dat_pre_data[751:744];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[93] | dat_pre_nan[46])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[751:744] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg7[759:752] <= dat_pre_data[759:752];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[94] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[759:752] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b1) begin
    dat_actv_data_reg7[767:760] <= dat_pre_data[767:760];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[95] | dat_pre_nan[47])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[767:760] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg7[775:768] <= dat_pre_data[775:768];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[96] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[775:768] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b1) begin
    dat_actv_data_reg7[783:776] <= dat_pre_data[783:776];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[97] | dat_pre_nan[48])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[783:776] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg7[791:784] <= dat_pre_data[791:784];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[98] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[791:784] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b1) begin
    dat_actv_data_reg7[799:792] <= dat_pre_data[799:792];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[99] | dat_pre_nan[49])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[799:792] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg7[807:800] <= dat_pre_data[807:800];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[100] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[807:800] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b1) begin
    dat_actv_data_reg7[815:808] <= dat_pre_data[815:808];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[101] | dat_pre_nan[50])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[815:808] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg7[823:816] <= dat_pre_data[823:816];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[102] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[823:816] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b1) begin
    dat_actv_data_reg7[831:824] <= dat_pre_data[831:824];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[103] | dat_pre_nan[51])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[831:824] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg7[839:832] <= dat_pre_data[839:832];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[104] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[839:832] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b1) begin
    dat_actv_data_reg7[847:840] <= dat_pre_data[847:840];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[105] | dat_pre_nan[52])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[847:840] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg7[855:848] <= dat_pre_data[855:848];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[106] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[855:848] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b1) begin
    dat_actv_data_reg7[863:856] <= dat_pre_data[863:856];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[107] | dat_pre_nan[53])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[863:856] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg7[871:864] <= dat_pre_data[871:864];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[108] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[871:864] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b1) begin
    dat_actv_data_reg7[879:872] <= dat_pre_data[879:872];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[109] | dat_pre_nan[54])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[879:872] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg7[887:880] <= dat_pre_data[887:880];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[110] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[887:880] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b1) begin
    dat_actv_data_reg7[895:888] <= dat_pre_data[895:888];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[111] | dat_pre_nan[55])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[895:888] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg7[903:896] <= dat_pre_data[903:896];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[112] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[903:896] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b1) begin
    dat_actv_data_reg7[911:904] <= dat_pre_data[911:904];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[113] | dat_pre_nan[56])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[911:904] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg7[919:912] <= dat_pre_data[919:912];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[114] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[919:912] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b1) begin
    dat_actv_data_reg7[927:920] <= dat_pre_data[927:920];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[115] | dat_pre_nan[57])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[927:920] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg7[935:928] <= dat_pre_data[935:928];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[116] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[935:928] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b1) begin
    dat_actv_data_reg7[943:936] <= dat_pre_data[943:936];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[117] | dat_pre_nan[58])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[943:936] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg7[951:944] <= dat_pre_data[951:944];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[118] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[951:944] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b1) begin
    dat_actv_data_reg7[959:952] <= dat_pre_data[959:952];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[119] | dat_pre_nan[59])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[959:952] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg7[967:960] <= dat_pre_data[967:960];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[120] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[967:960] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b1) begin
    dat_actv_data_reg7[975:968] <= dat_pre_data[975:968];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[121] | dat_pre_nan[60])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[975:968] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg7[983:976] <= dat_pre_data[983:976];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[122] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[983:976] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b1) begin
    dat_actv_data_reg7[991:984] <= dat_pre_data[991:984];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[123] | dat_pre_nan[61])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[991:984] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg7[999:992] <= dat_pre_data[999:992];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[124] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[999:992] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b1) begin
    dat_actv_data_reg7[1007:1000] <= dat_pre_data[1007:1000];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[125] | dat_pre_nan[62])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[1007:1000] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg7[1015:1008] <= dat_pre_data[1015:1008];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[126] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[1015:1008] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end
always @(posedge nvdla_core_clk) begin
  if ((dat_pre_pvld[15] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b1) begin
    dat_actv_data_reg7[1023:1016] <= dat_pre_data[1023:1016];
  // VCS coverage off
  end else if ((dat_pre_pvld[15] & (dat_pre_nz[127] | dat_pre_nan[63])) == 1'b0) begin
  end else begin
    dat_actv_data_reg7[1023:1016] <= 'bx;  // spyglass disable STARC-2.10.1.6 W443 NoWidthInBasedNum-ML -- (Constant containing x or z used, Based number `bx contains an X, Width specification missing for based number)
  // VCS coverage on
  end
end










always @(
  dat_actv_pvld_reg0
  or dat_actv_data_reg0
  or dat_actv_nz_reg0
  or dat_actv_nan_reg0
  ) begin
    dat0_actv_pvld = dat_actv_pvld_reg0;
    dat0_actv_data = dat_actv_data_reg0;
    dat0_actv_nz   = dat_actv_nz_reg0;
    dat0_actv_nan  = dat_actv_nan_reg0;
end




always @(
  dat_actv_pvld_reg1
  or dat_actv_data_reg1
  or dat_actv_nz_reg1
  or dat_actv_nan_reg1
  ) begin
    dat1_actv_pvld = dat_actv_pvld_reg1;
    dat1_actv_data = dat_actv_data_reg1;
    dat1_actv_nz   = dat_actv_nz_reg1;
    dat1_actv_nan  = dat_actv_nan_reg1;
end




always @(
  dat_actv_pvld_reg2
  or dat_actv_data_reg2
  or dat_actv_nz_reg2
  or dat_actv_nan_reg2
  ) begin
    dat2_actv_pvld = dat_actv_pvld_reg2;
    dat2_actv_data = dat_actv_data_reg2;
    dat2_actv_nz   = dat_actv_nz_reg2;
    dat2_actv_nan  = dat_actv_nan_reg2;
end




always @(
  dat_actv_pvld_reg3
  or dat_actv_data_reg3
  or dat_actv_nz_reg3
  or dat_actv_nan_reg3
  ) begin
    dat3_actv_pvld = dat_actv_pvld_reg3;
    dat3_actv_data = dat_actv_data_reg3;
    dat3_actv_nz   = dat_actv_nz_reg3;
    dat3_actv_nan  = dat_actv_nan_reg3;
end




always @(
  dat_actv_pvld_reg4
  or dat_actv_data_reg4
  or dat_actv_nz_reg4
  or dat_actv_nan_reg4
  ) begin
    dat4_actv_pvld = dat_actv_pvld_reg4;
    dat4_actv_data = dat_actv_data_reg4;
    dat4_actv_nz   = dat_actv_nz_reg4;
    dat4_actv_nan  = dat_actv_nan_reg4;
end




always @(
  dat_actv_pvld_reg5
  or dat_actv_data_reg5
  or dat_actv_nz_reg5
  or dat_actv_nan_reg5
  ) begin
    dat5_actv_pvld = dat_actv_pvld_reg5;
    dat5_actv_data = dat_actv_data_reg5;
    dat5_actv_nz   = dat_actv_nz_reg5;
    dat5_actv_nan  = dat_actv_nan_reg5;
end




always @(
  dat_actv_pvld_reg6
  or dat_actv_data_reg6
  or dat_actv_nz_reg6
  or dat_actv_nan_reg6
  ) begin
    dat6_actv_pvld = dat_actv_pvld_reg6;
    dat6_actv_data = dat_actv_data_reg6;
    dat6_actv_nz   = dat_actv_nz_reg6;
    dat6_actv_nan  = dat_actv_nan_reg6;
end




always @(
  dat_actv_pvld_reg7
  or dat_actv_data_reg7
  or dat_actv_nz_reg7
  or dat_actv_nan_reg7
  ) begin
    dat7_actv_pvld = dat_actv_pvld_reg7;
    dat7_actv_data = dat_actv_data_reg7;
    dat7_actv_nz   = dat_actv_nz_reg7;
    dat7_actv_nan  = dat_actv_nan_reg7;
end




endmodule // NV_NVDLA_CMAC_CORE_active


