// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: HLS_fp17_mul.v

module FP17_MUL_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/FP17_MUL_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module FP17_MUL_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-184
//  Generated date: Fri Jun 16 21:52:26 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP17_MUL_chn_o_rsci_unreg
// ------------------------------------------------------------------


module FP17_MUL_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP17_MUL_chn_b_rsci_unreg
// ------------------------------------------------------------------


module FP17_MUL_chn_b_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP17_MUL_chn_a_rsci_unreg
// ------------------------------------------------------------------


module FP17_MUL_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module HLS_fp17_mul_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for HLS_fp17_mul_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : HLS_fp17_mul_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_staller
// ------------------------------------------------------------------


module HLS_fp17_mul_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_b_rsci_wen_comp,
      chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_b_rsci_wen_comp;
  input chn_o_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_a_rsci_wen_comp & chn_b_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;


  // Interconnect Declarations
  reg chn_o_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;


  // Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_d_mxwt, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  output [16:0] chn_b_rsci_d_mxwt;
  input chn_b_rsci_biwt;
  input chn_b_rsci_bdwt;
  input [16:0] chn_b_rsci_d;


  // Interconnect Declarations
  reg chn_b_rsci_bcwt;
  reg [16:0] chn_b_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_bawt = chn_b_rsci_biwt | chn_b_rsci_bcwt;
  assign chn_b_rsci_wen_comp = (~ chn_b_rsci_oswt) | chn_b_rsci_bawt;
  assign chn_b_rsci_d_mxwt = MUX_v_17_2_2(chn_b_rsci_d, chn_b_rsci_d_bfwt, chn_b_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_bcwt <= 1'b0;
      chn_b_rsci_d_bfwt <= 17'b0;
    end
    else begin
      chn_b_rsci_bcwt <= ~((~(chn_b_rsci_bcwt | chn_b_rsci_biwt)) | chn_b_rsci_bdwt);
      chn_b_rsci_d_bfwt <= chn_b_rsci_d_mxwt;
    end
  end

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, core_wen, core_wten, chn_b_rsci_iswt0,
      chn_b_rsci_ld_core_psct, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_ld_core_sct,
      chn_b_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  input chn_b_rsci_ld_core_psct;
  output chn_b_rsci_biwt;
  output chn_b_rsci_bdwt;
  output chn_b_rsci_ld_core_sct;
  input chn_b_rsci_vd;


  // Interconnect Declarations
  wire chn_b_rsci_ogwt;
  wire chn_b_rsci_pdswt0;
  reg chn_b_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_pdswt0 = (~ core_wten) & chn_b_rsci_iswt0;
  assign chn_b_rsci_biwt = chn_b_rsci_ogwt & chn_b_rsci_vd;
  assign chn_b_rsci_ogwt = chn_b_rsci_pdswt0 | chn_b_rsci_icwt;
  assign chn_b_rsci_bdwt = chn_b_rsci_oswt & core_wen;
  assign chn_b_rsci_ld_core_sct = chn_b_rsci_ld_core_psct & chn_b_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_icwt <= 1'b0;
    end
    else begin
      chn_b_rsci_icwt <= ~((~(chn_b_rsci_icwt | chn_b_rsci_pdswt0)) | chn_b_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [16:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [16:0] chn_a_rsci_d;


  // Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [16:0] chn_a_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_17_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 17'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;


  // Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_o_rsci
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [16:0] chn_o_rsci_d;


  // Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  FP17_MUL_mgc_out_stdreg_wait_v1 #(.rscid(32'sd3),
  .width(32'sd17)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(chn_o_rsci_d),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_ctrl HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_dp HLS_fp17_mul_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_b_rsci
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_b_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsc_z, chn_b_rsc_vz, chn_b_rsc_lz, chn_b_rsci_oswt,
      core_wen, core_wten, chn_b_rsci_iswt0, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_ld_core_psct, chn_b_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  input chn_b_rsci_ld_core_psct;
  output [16:0] chn_b_rsci_d_mxwt;


  // Interconnect Declarations
  wire chn_b_rsci_biwt;
  wire chn_b_rsci_bdwt;
  wire chn_b_rsci_ld_core_sct;
  wire chn_b_rsci_vd;
  wire [16:0] chn_b_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP17_MUL_mgc_in_wire_wait_v1 #(.rscid(32'sd2),
  .width(32'sd17)) chn_b_rsci (
      .ld(chn_b_rsci_ld_core_sct),
      .vd(chn_b_rsci_vd),
      .d(chn_b_rsci_d),
      .lz(chn_b_rsc_lz),
      .vz(chn_b_rsc_vz),
      .z(chn_b_rsc_z)
    );
  HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_ctrl HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(chn_b_rsci_iswt0),
      .chn_b_rsci_ld_core_psct(chn_b_rsci_ld_core_psct),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_ld_core_sct(chn_b_rsci_ld_core_sct),
      .chn_b_rsci_vd(chn_b_rsci_vd)
    );
  HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_dp HLS_fp17_mul_core_chn_b_rsci_chn_b_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_d(chn_b_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core_chn_a_rsci
// ------------------------------------------------------------------


module HLS_fp17_mul_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [16:0] chn_a_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [16:0] chn_a_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP17_MUL_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd17)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_ctrl HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_dp HLS_fp17_mul_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul_core
// ------------------------------------------------------------------


module HLS_fp17_mul_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt,
      chn_b_rsci_oswt, chn_o_rsci_oswt, chn_o_rsci_oswt_unreg, chn_a_rsci_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  input chn_b_rsci_oswt;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;
  output chn_a_rsci_oswt_unreg_pff;


  // Interconnect Declarations
  wire core_wen;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  wire [16:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  wire chn_b_rsci_bawt;
  wire chn_b_rsci_wen_comp;
  wire [16:0] chn_b_rsci_d_mxwt;
  reg chn_o_rsci_iswt0;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg chn_o_rsci_d_16;
  reg [5:0] chn_o_rsci_d_15_10;
  reg [9:0] chn_o_rsci_d_9_0;
  wire [1:0] fsm_output;
  wire IsNaN_6U_10U_nor_tmp;
  wire FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp;
  wire [21:0] FpMul_6U_10U_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_1_nor_tmp;
  wire nor_tmp_1;
  wire or_tmp_4;
  wire mux_tmp_3;
  wire or_tmp_7;
  wire or_tmp_16;
  wire mux_tmp_6;
  wire mux_tmp_7;
  wire nor_tmp_11;
  wire or_tmp_32;
  wire or_tmp_40;
  wire mux_tmp_21;
  wire mux_tmp_23;
  wire or_tmp_48;
  wire or_tmp_49;
  wire or_tmp_52;
  wire and_dcpl_7;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_28;
  wire or_tmp_56;
  wire or_tmp_62;
  wire or_tmp_68;
  reg FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_p_mant_p1_sva;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_3;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_4;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_3;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_4;
  reg FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_3;
  reg FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_4;
  reg [21:0] FpMul_6U_10U_p_mant_p1_sva_2;
  reg [5:0] FpMul_6U_10U_p_expo_sva_5;
  wire [6:0] nl_FpMul_6U_10U_p_expo_sva_5;
  reg IsNaN_6U_10U_land_lpi_1_dfm_4;
  reg [5:0] FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_15_10_itm_2;
  reg FpMul_6U_10U_mux_10_itm_3;
  reg FpMul_6U_10U_mux_10_itm_4;
  reg [9:0] FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_9_0_itm_2;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_st_4;
  reg FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4;
  reg FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2;
  reg IsNaN_6U_10U_land_lpi_1_dfm_st_3;
  reg [15:0] FpMul_6U_10U_ua_sva_1_15_0_1;
  reg [15:0] FpMul_6U_10U_ub_sva_1_15_0_1;
  wire main_stage_en_1;
  wire FpMantRNE_22U_11U_else_and_svs;
  wire FpMul_6U_10U_is_inf_lpi_1_dfm_2;
  wire FpMantRNE_22U_11U_else_carry_sva;
  wire [5:0] FpMul_6U_10U_o_expo_lpi_1_dfm;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1;
  wire [19:0] FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0;
  reg reg_chn_b_rsci_iswt0_cse;
  reg reg_chn_b_rsci_ld_core_psct_cse;
  wire chn_o_and_cse;
  wire nor_42_cse;
  wire or_65_cse;
  wire nor_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire or_68_cse;
  wire or_5_cse;
  wire nand_cse;
  wire FpMul_6U_10U_or_2_cse;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_nand_cse;
  wire nand_7_cse;
  wire nand_6_cse;
  wire and_40_rgt;
  wire and_45_rgt;
  wire and_52_rgt;
  wire and_60_rgt;
  wire and_61_rgt;
  wire chn_o_rsci_d_15_10_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire [5:0] FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0;
  wire FpMul_6U_10U_lor_2_lpi_1_dfm;
  wire IsNaN_6U_10U_aelse_and_cse;
  wire IsNaN_6U_10U_1_aelse_and_cse;
  wire FpMul_6U_10U_oelse_1_and_1_cse;
  wire FpBitsToFloat_6U_10U_1_and_1_cse;
  wire FpMul_6U_10U_else_2_if_acc_itm_6_1;
  wire FpMul_6U_10U_oelse_1_acc_itm_7_1;
  wire FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1;

  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[9:0] FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_1_nl;
  wire[9:0] FpMul_6U_10U_nor_nl;
  wire[9:0] mux_37_nl;
  wire[9:0] FpMantRNE_22U_11U_else_acc_nl;
  wire[10:0] nl_FpMantRNE_22U_11U_else_acc_nl;
  wire[0:0] or_nl;
  wire[5:0] FpMul_6U_10U_FpMul_6U_10U_and_2_nl;
  wire[0:0] FpMul_6U_10U_oelse_2_not_1_nl;
  wire[0:0] FpBitsToFloat_6U_10U_1_and_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] or_2_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] mux_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_acc_2_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_acc_2_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_41_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_43_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] nor_39_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] nor_38_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] nor_6_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_25_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] nor_37_nl;
  wire[0:0] and_97_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] or_35_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] or_38_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] and_91_nl;
  wire[0:0] FpMul_6U_10U_xor_1_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] nor_33_nl;
  wire[6:0] FpMul_6U_10U_else_2_if_acc_nl;
  wire[7:0] nl_FpMul_6U_10U_else_2_if_acc_nl;
  wire[6:0] FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] nl_FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] FpMul_6U_10U_oelse_1_acc_nl;
  wire[8:0] nl_FpMul_6U_10U_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_oelse_1_acc_1_nl;
  wire[7:0] nl_FpMul_6U_10U_oelse_1_acc_1_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[0:0] and_62_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_nor_1_nl;
  wire[0:0] FpMul_6U_10U_or_1_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] and_93_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] and_94_nl;
  wire[0:0] nor_34_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [16:0] nl_HLS_fp17_mul_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_fp17_mul_core_chn_o_rsci_inst_chn_o_rsci_d = {chn_o_rsci_d_16 , chn_o_rsci_d_15_10
      , chn_o_rsci_d_9_0};
  HLS_fp17_mul_core_chn_a_rsci HLS_fp17_mul_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_fp17_mul_core_chn_b_rsci HLS_fp17_mul_core_chn_b_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt)
    );
  HLS_fp17_mul_core_chn_o_rsci HLS_fp17_mul_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_fp17_mul_core_chn_o_rsci_inst_chn_o_rsci_d[16:0])
    );
  HLS_fp17_mul_core_staller HLS_fp17_mul_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_fp17_mul_core_core_fsm HLS_fp17_mul_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign iMantWidth_oMantWidth_prb = MUX_s_1_2_2((MUX1HOT_s_1_1_2(1'b1, fsm_output[0])),
      (MUX1HOT_s_1_1_2(1'b1, main_stage_en_1 & (fsm_output[1]))), fsm_output[1]);
  // assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 386
  // PSL HLS_fp17_mul_core_nvdla_float_h_ln386_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign chn_o_and_cse = core_wen & (~(and_dcpl_7 | (~ main_stage_v_2)));
  assign FpMul_6U_10U_or_2_cse = IsNaN_6U_10U_1_land_lpi_1_dfm_4 | IsNaN_6U_10U_land_lpi_1_dfm_4;
  assign nor_cse = ~(chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign IsNaN_6U_10U_aelse_and_cse = core_wen & (~ and_dcpl_7) & mux_tmp_3;
  assign nor_42_cse = ~((~ main_stage_v_2) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 |
      (~ FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4));
  assign or_5_cse = (~ reg_chn_o_rsci_ld_core_psct_cse) | chn_o_rsci_bawt;
  assign or_65_cse = FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 | (~ FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3);
  assign and_40_rgt = or_5_cse & or_65_cse;
  assign or_25_nl = nor_cse | nor_tmp_11;
  assign nor_37_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ nor_tmp_11));
  assign mux_12_nl = MUX_s_1_2_2((nor_37_nl), nor_tmp_11, chn_o_rsci_bawt);
  assign and_97_nl = FpMul_6U_10U_or_2_cse & main_stage_v_2;
  assign mux_13_nl = MUX_s_1_2_2((mux_12_nl), (or_25_nl), and_97_nl);
  assign FpBitsToFloat_6U_10U_1_and_1_cse = core_wen & ((or_5_cse & (~ IsNaN_6U_10U_land_lpi_1_dfm_st_3))
      | and_dcpl_28) & (mux_13_nl);
  assign IsNaN_6U_10U_1_aelse_and_cse = core_wen & (~ and_dcpl_7) & mux_tmp_7;
  assign nor_35_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ or_tmp_32));
  assign mux_16_nl = MUX_s_1_2_2((nor_35_nl), or_tmp_32, chn_o_rsci_bawt);
  assign or_35_nl = nor_cse | IsNaN_6U_10U_1_land_lpi_1_dfm_3 | IsNaN_6U_10U_land_lpi_1_dfm_st_3
      | (~ main_stage_v_1);
  assign nor_15_nl = ~(IsNaN_6U_10U_1_land_lpi_1_dfm_4 | IsNaN_6U_10U_land_lpi_1_dfm_4
      | (~ main_stage_v_2));
  assign mux_17_nl = MUX_s_1_2_2((or_35_nl), (mux_16_nl), nor_15_nl);
  assign FpMul_6U_10U_oelse_1_and_1_cse = core_wen & (~ and_dcpl_7) & (~ (mux_17_nl));
  assign or_68_cse = FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp | FpMul_6U_10U_oelse_1_acc_itm_7_1;
  assign and_45_rgt = or_68_cse & or_5_cse;
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_nand_cse = ~((chn_b_rsci_d_mxwt[15:10]==6'b111111));
  assign nand_cse = ~((chn_a_rsci_d_mxwt[15:10]==6'b111111));
  assign and_52_rgt = or_5_cse & (chn_a_rsci_d_mxwt[15:10]==6'b111111) & (~ IsNaN_6U_10U_nor_tmp);
  assign and_60_rgt = ((chn_a_rsci_d_mxwt[15:10]!=6'b111111) | IsNaN_6U_10U_nor_tmp)
      & (chn_b_rsci_d_mxwt[15:10]==6'b111111) & (~ IsNaN_6U_10U_1_nor_tmp) & or_5_cse;
  assign and_91_nl = nand_cse & or_tmp_56;
  assign mux_35_nl = MUX_s_1_2_2((and_91_nl), or_tmp_56, IsNaN_6U_10U_nor_tmp);
  assign and_61_rgt = (mux_35_nl) & or_5_cse;
  assign nand_7_cse = ~(FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3
      & main_stage_v_1);
  assign nand_6_cse = ~(chn_a_rsci_bawt & chn_b_rsci_bawt);
  assign nl_FpMul_6U_10U_else_2_acc_1_nl = conv_u2u_6_7(chn_a_rsci_d_mxwt[15:10])
      + conv_u2u_6_7(chn_b_rsci_d_mxwt[15:10]);
  assign FpMul_6U_10U_else_2_acc_1_nl = nl_FpMul_6U_10U_else_2_acc_1_nl[6:0];
  assign nl_FpMul_6U_10U_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((FpMul_6U_10U_else_2_acc_1_nl)))
      + 7'b1010001;
  assign FpMul_6U_10U_else_2_if_acc_nl = nl_FpMul_6U_10U_else_2_if_acc_nl[6:0];
  assign FpMul_6U_10U_else_2_if_acc_itm_6_1 = readslicef_7_1_6((FpMul_6U_10U_else_2_if_acc_nl));
  assign IsNaN_6U_10U_nor_tmp = ~((chn_a_rsci_d_mxwt[9:0]!=10'b0000000000));
  assign FpMul_6U_10U_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 , (FpMul_6U_10U_ua_sva_1_15_0_1[9:0])})
      * ({1'b1 , (FpMul_6U_10U_ub_sva_1_15_0_1[9:0])}));
  assign IsNaN_6U_10U_1_nor_tmp = ~((chn_b_rsci_d_mxwt[9:0]!=10'b0000000000));
  assign nl_FpMul_6U_10U_oelse_1_acc_1_nl = conv_u2s_6_7(chn_b_rsci_d_mxwt[15:10])
      + 7'b1100001;
  assign FpMul_6U_10U_oelse_1_acc_1_nl = nl_FpMul_6U_10U_oelse_1_acc_1_nl[6:0];
  assign nl_FpMul_6U_10U_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_oelse_1_acc_1_nl)
      + conv_u2s_6_8(chn_a_rsci_d_mxwt[15:10]);
  assign FpMul_6U_10U_oelse_1_acc_nl = nl_FpMul_6U_10U_oelse_1_acc_nl[7:0];
  assign FpMul_6U_10U_oelse_1_acc_itm_7_1 = readslicef_8_1_7((FpMul_6U_10U_oelse_1_acc_nl));
  assign FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp = (~((chn_b_rsci_d_mxwt[15:0]!=16'b0000000000000000)))
      | (~((chn_a_rsci_d_mxwt[15:0]!=16'b0000000000000000)));
  assign nl_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_p_expo_sva_5[5:1])})
      + 6'b1;
  assign FpMul_6U_10U_else_2_else_if_if_acc_1_nl = nl_FpMul_6U_10U_else_2_else_if_if_acc_1_nl[5:0];
  assign FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((FpMul_6U_10U_else_2_else_if_if_acc_1_nl));
  assign nl_FpMul_6U_10U_else_2_else_if_if_acc_nl = FpMul_6U_10U_p_expo_sva_5 + 6'b1;
  assign FpMul_6U_10U_else_2_else_if_if_acc_nl = nl_FpMul_6U_10U_else_2_else_if_if_acc_nl[5:0];
  assign mux_36_nl = MUX_s_1_2_2((~ FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2),
      FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2, FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1);
  assign and_62_nl = (mux_36_nl) & (FpMul_6U_10U_p_mant_p1_sva_2[21]);
  assign FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(FpMul_6U_10U_p_expo_sva_5,
      (FpMul_6U_10U_else_2_else_if_if_acc_nl), and_62_nl);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp = ~((FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1 = FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1[5:0];
  assign FpMantRNE_22U_11U_else_and_svs = FpMantRNE_22U_11U_else_carry_sva & (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMantRNE_22U_11U_else_carry_sva = (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_p_mant_p1_sva_2[0]) & (FpMul_6U_10U_p_mant_p1_sva_2[21]))
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[10]));
  assign FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_p_mant_p1_sva_2[19:0]),
      (FpMul_6U_10U_p_mant_p1_sva_2[20:1]), FpMul_6U_10U_p_mant_p1_sva_2[21]);
  assign FpMul_6U_10U_FpMul_6U_10U_nor_1_nl = ~(FpMantRNE_22U_11U_else_and_svs |
      FpMul_6U_10U_is_inf_lpi_1_dfm_2);
  assign FpMul_6U_10U_or_1_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp)
      & FpMantRNE_22U_11U_else_and_svs) | FpMul_6U_10U_is_inf_lpi_1_dfm_2;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp
      & FpMantRNE_22U_11U_else_and_svs & (~ FpMul_6U_10U_is_inf_lpi_1_dfm_2);
  assign FpMul_6U_10U_o_expo_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1, {(FpMul_6U_10U_FpMul_6U_10U_nor_1_nl)
      , (FpMul_6U_10U_or_1_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl)});
  assign FpMul_6U_10U_lor_2_lpi_1_dfm = (~((FpMul_6U_10U_o_expo_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_lor_1_lpi_1_dfm_4;
  assign FpMul_6U_10U_is_inf_lpi_1_dfm_2 = ~(((FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      | (~ (FpMul_6U_10U_p_mant_p1_sva_2[21]))) & FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_4)
      | FpMul_6U_10U_lor_1_lpi_1_dfm_4);
  assign main_stage_en_1 = chn_a_rsci_bawt & chn_b_rsci_bawt & or_5_cse;
  assign nor_tmp_1 = chn_a_rsci_bawt & chn_b_rsci_bawt;
  assign or_tmp_4 = FpMul_6U_10U_oelse_1_acc_itm_7_1 | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp
      | (~ nor_tmp_1);
  assign mux_tmp_3 = MUX_s_1_2_2(nor_tmp_1, main_stage_v_1, nor_cse);
  assign or_tmp_7 = IsNaN_6U_10U_land_lpi_1_dfm_st_3 | IsNaN_6U_10U_1_land_lpi_1_dfm_3;
  assign or_tmp_16 = nor_cse | main_stage_v_1;
  assign nor_40_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ main_stage_v_1));
  assign mux_tmp_6 = MUX_s_1_2_2((nor_40_nl), main_stage_v_1, chn_o_rsci_bawt);
  assign mux_tmp_7 = MUX_s_1_2_2(mux_tmp_6, or_tmp_16, main_stage_v_2);
  assign nor_tmp_11 = or_tmp_7 & main_stage_v_1;
  assign or_tmp_32 = or_tmp_7 | (~ main_stage_v_1);
  assign or_tmp_40 = (~ FpMul_6U_10U_else_2_if_acc_itm_6_1) | FpMul_6U_10U_oelse_1_acc_itm_7_1
      | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp | (~ nor_tmp_1);
  assign and_93_nl = nand_cse & nor_tmp_1;
  assign mux_tmp_21 = MUX_s_1_2_2((and_93_nl), nor_tmp_1, IsNaN_6U_10U_nor_tmp);
  assign and_94_nl = IsNaN_6U_10U_1_IsNaN_6U_10U_1_nand_cse & mux_tmp_21;
  assign mux_22_nl = MUX_s_1_2_2((and_94_nl), mux_tmp_21, IsNaN_6U_10U_1_nor_tmp);
  assign nor_34_nl = ~((~ main_stage_v_1) | IsNaN_6U_10U_land_lpi_1_dfm_st_3 | IsNaN_6U_10U_1_land_lpi_1_dfm_3);
  assign mux_tmp_23 = MUX_s_1_2_2((nor_34_nl), (mux_22_nl), or_5_cse);
  assign or_tmp_48 = IsNaN_6U_10U_1_nor_tmp | (~((chn_b_rsci_d_mxwt[15:10]==6'b111111)
      & mux_tmp_21));
  assign or_tmp_49 = FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 | nand_7_cse;
  assign or_tmp_52 = IsNaN_6U_10U_nor_tmp | (~((chn_a_rsci_d_mxwt[15:10]==6'b111111)
      & chn_a_rsci_bawt & chn_b_rsci_bawt));
  assign and_dcpl_7 = reg_chn_o_rsci_ld_core_psct_cse & (~ chn_o_rsci_bawt);
  assign and_dcpl_13 = or_5_cse & main_stage_v_2;
  assign and_dcpl_14 = reg_chn_o_rsci_ld_core_psct_cse & chn_o_rsci_bawt;
  assign and_dcpl_15 = and_dcpl_14 & (~ main_stage_v_2);
  assign and_dcpl_28 = or_5_cse & IsNaN_6U_10U_land_lpi_1_dfm_st_3;
  assign or_tmp_56 = IsNaN_6U_10U_1_nor_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_nand_cse;
  assign or_tmp_62 = main_stage_en_1 | (fsm_output[0]);
  assign or_tmp_68 = chn_b_rsci_bawt & chn_a_rsci_bawt & or_5_cse & (fsm_output[1]);
  assign chn_o_rsci_d_15_10_mx0c1 = or_5_cse & main_stage_v_2 & (~ IsNaN_6U_10U_land_lpi_1_dfm_4);
  assign main_stage_v_1_mx0c1 = nand_6_cse & main_stage_v_1 & or_5_cse;
  assign main_stage_v_2_mx0c1 = or_5_cse & (~ main_stage_v_1) & main_stage_v_2;
  assign chn_a_rsci_oswt_unreg_pff = or_tmp_68;
  assign chn_o_rsci_oswt_unreg = and_dcpl_14;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_iswt0_cse <= 1'b0;
      chn_o_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_chn_b_rsci_iswt0_cse <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_o_rsci_iswt0 <= and_dcpl_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & or_tmp_62 ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= or_tmp_62;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_9_0 <= 10'b0;
      chn_o_rsci_d_16 <= 1'b0;
    end
    else if ( chn_o_and_cse ) begin
      chn_o_rsci_d_9_0 <= MUX_v_10_2_2((FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_1_nl),
          FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_9_0_itm_2, FpMul_6U_10U_or_2_cse);
      chn_o_rsci_d_16 <= FpMul_6U_10U_mux_10_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_15_10 <= 6'b0;
    end
    else if ( core_wen & ((or_5_cse & main_stage_v_2 & IsNaN_6U_10U_land_lpi_1_dfm_4)
        | chn_o_rsci_d_15_10_mx0c1) ) begin
      chn_o_rsci_d_15_10 <= MUX_v_6_2_2(FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_15_10_itm_2,
          (FpMul_6U_10U_FpMul_6U_10U_and_2_nl), FpBitsToFloat_6U_10U_1_and_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_13 | and_dcpl_15) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_68 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (~ (mux_2_nl)) ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3 <= FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_land_lpi_1_dfm_st_3 <= 1'b0;
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_1_land_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_aelse_and_cse ) begin
      IsNaN_6U_10U_land_lpi_1_dfm_st_3 <= ~(IsNaN_6U_10U_nor_tmp | nand_cse);
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 <= or_68_cse;
      IsNaN_6U_10U_1_land_lpi_1_dfm_3 <= ~(IsNaN_6U_10U_1_nor_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_nand_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5_cse & main_stage_v_1) | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_expo_sva_5 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_5_nl) ) begin
      FpMul_6U_10U_p_expo_sva_5 <= nl_FpMul_6U_10U_p_expo_sva_5[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_sva_2 <= 22'b0;
    end
    else if ( core_wen & ((or_5_cse & (~ FpMul_6U_10U_lor_1_lpi_1_dfm_st_3) & FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3)
        | and_40_rgt) & mux_tmp_7 ) begin
      FpMul_6U_10U_p_mant_p1_sva_2 <= MUX_v_22_2_2(FpMul_6U_10U_p_mant_p1_mul_tmp,
          FpMul_6U_10U_p_mant_p1_sva, and_40_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_9_nl) ) begin
      FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <= FpMul_6U_10U_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_11_nl) ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4 <= FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_15_10_itm_2 <= 6'b0;
      FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_9_0_itm_2 <= 10'b0;
    end
    else if ( FpBitsToFloat_6U_10U_1_and_1_cse ) begin
      FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_15_10_itm_2 <= MUX_v_6_2_2((FpMul_6U_10U_ub_sva_1_15_0_1[15:10]),
          (FpMul_6U_10U_ua_sva_1_15_0_1[15:10]), and_dcpl_28);
      FpBitsToFloat_6U_10U_1_slc_FpBitsToFloat_6U_10U_ubits_1_9_0_itm_2 <= MUX_v_10_2_2((FpMul_6U_10U_ub_sva_1_15_0_1[9:0]),
          (FpMul_6U_10U_ua_sva_1_15_0_1[9:0]), and_dcpl_28);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_4 <= 1'b0;
      FpMul_6U_10U_mux_10_itm_4 <= 1'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_4 <= 1'b0;
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_1_aelse_and_cse ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_4 <= IsNaN_6U_10U_1_land_lpi_1_dfm_3;
      FpMul_6U_10U_mux_10_itm_4 <= FpMul_6U_10U_mux_10_itm_3;
      IsNaN_6U_10U_land_lpi_1_dfm_4 <= IsNaN_6U_10U_land_lpi_1_dfm_st_3;
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 <= FpMul_6U_10U_lor_1_lpi_1_dfm_st_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_4 <= 1'b0;
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_4 <= 1'b0;
    end
    else if ( FpMul_6U_10U_oelse_1_and_1_cse ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_4 <= FpMul_6U_10U_lor_1_lpi_1_dfm_3;
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_4 <= FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_sva <= 22'b0;
    end
    else if ( core_wen & (~ (fsm_output[0])) & (~((~ main_stage_v_1) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_3
        | (~ FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3)))
        & (mux_20_nl) ) begin
      FpMul_6U_10U_p_mant_p1_sva <= FpMul_6U_10U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & mux_tmp_23 ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_3 <= or_68_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_3 <= 1'b0;
    end
    else if ( core_wen & (((~(FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp | FpMul_6U_10U_oelse_1_acc_itm_7_1))
        & or_5_cse) | and_45_rgt) & mux_tmp_23 ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_3 <= MUX_s_1_2_2(FpMul_6U_10U_else_2_if_acc_itm_6_1,
          FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs, and_45_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_mux_10_itm_3 <= 1'b0;
    end
    else if ( core_wen & (and_52_rgt | and_60_rgt | and_61_rgt) & mux_tmp_3 ) begin
      FpMul_6U_10U_mux_10_itm_3 <= MUX1HOT_s_1_3_2((chn_a_rsci_d_mxwt[16]), (chn_b_rsci_d_mxwt[16]),
          (FpMul_6U_10U_xor_1_nl), {and_52_rgt , and_60_rgt , and_61_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_ub_sva_1_15_0_1 <= 16'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (~ (mux_29_nl)) ) begin
      FpMul_6U_10U_ub_sva_1_15_0_1 <= chn_b_rsci_d_mxwt[15:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_ua_sva_1_15_0_1 <= 16'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_33_nl) ) begin
      FpMul_6U_10U_ua_sva_1_15_0_1 <= chn_a_rsci_d_mxwt[15:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <= 1'b0;
    end
    else if ( core_wen & (~(nand_6_cse | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp
        | and_dcpl_7 | FpMul_6U_10U_oelse_1_acc_itm_7_1 | (fsm_output[0]))) ) begin
      FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <= FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  assign nl_FpMantRNE_22U_11U_else_acc_nl = (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[19:10])
      + conv_u2u_1_10(FpMantRNE_22U_11U_else_carry_sva);
  assign FpMantRNE_22U_11U_else_acc_nl = nl_FpMantRNE_22U_11U_else_acc_nl[9:0];
  assign or_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp | (~ FpMantRNE_22U_11U_else_and_svs);
  assign mux_37_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp)),
      (FpMantRNE_22U_11U_else_acc_nl), or_nl);
  assign FpMul_6U_10U_nor_nl = ~(MUX_v_10_2_2((mux_37_nl), 10'b1111111111, FpMul_6U_10U_is_inf_lpi_1_dfm_2));
  assign FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_1_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_nor_nl),
      10'b1111111111, FpMul_6U_10U_lor_2_lpi_1_dfm));
  assign FpMul_6U_10U_oelse_2_not_1_nl = ~ FpMul_6U_10U_lor_2_lpi_1_dfm;
  assign FpMul_6U_10U_FpMul_6U_10U_and_2_nl = MUX_v_6_2_2(6'b000000, FpMul_6U_10U_o_expo_lpi_1_dfm,
      (FpMul_6U_10U_oelse_2_not_1_nl));
  assign FpBitsToFloat_6U_10U_1_and_nl = (~ IsNaN_6U_10U_1_land_lpi_1_dfm_4) & chn_o_rsci_d_15_10_mx0c1;
  assign or_2_nl = nor_cse | FpMul_6U_10U_oelse_1_acc_itm_7_1 | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp
      | (~ nor_tmp_1);
  assign mux_nl = MUX_s_1_2_2(or_tmp_4, (~ main_stage_v_1), reg_chn_o_rsci_ld_core_psct_cse);
  assign mux_1_nl = MUX_s_1_2_2((mux_nl), or_tmp_4, chn_o_rsci_bawt);
  assign mux_2_nl = MUX_s_1_2_2((mux_1_nl), (or_2_nl), FpMul_6U_10U_lor_1_lpi_1_dfm_st_3);
  assign nl_FpMul_6U_10U_else_2_else_acc_2_nl = (FpMul_6U_10U_ub_sva_1_15_0_1[15:10])
      + 6'b100001;
  assign FpMul_6U_10U_else_2_else_acc_2_nl = nl_FpMul_6U_10U_else_2_else_acc_2_nl[5:0];
  assign nl_FpMul_6U_10U_p_expo_sva_5  = (FpMul_6U_10U_else_2_else_acc_2_nl) + (FpMul_6U_10U_ua_sva_1_15_0_1[15:10]);
  assign nor_41_nl = ~((~ main_stage_v_1) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 | (~(FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_3
      & ((FpMul_6U_10U_p_mant_p1_mul_tmp[21]) | (~ or_tmp_7)))));
  assign nor_43_nl = ~(FpMul_6U_10U_or_2_cse | (FpMul_6U_10U_p_mant_p1_sva_2[21])
      | (~ main_stage_v_2) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 | (~ FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4));
  assign mux_4_nl = MUX_s_1_2_2((nor_43_nl), nor_42_cse, FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2);
  assign mux_5_nl = MUX_s_1_2_2((mux_4_nl), (nor_41_nl), or_5_cse);
  assign nor_39_nl = ~((~ FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 | (~ main_stage_v_2) | chn_o_rsci_bawt
      | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign mux_8_nl = MUX_s_1_2_2(mux_tmp_6, or_tmp_16, nor_42_cse);
  assign mux_9_nl = MUX_s_1_2_2((mux_8_nl), (nor_39_nl), or_65_cse);
  assign nor_38_nl = ~(FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 | (~ main_stage_v_2) | chn_o_rsci_bawt
      | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign nor_6_nl = ~(FpMul_6U_10U_lor_1_lpi_1_dfm_st_4 | (~ main_stage_v_2));
  assign mux_10_nl = MUX_s_1_2_2(mux_tmp_6, or_tmp_16, nor_6_nl);
  assign mux_11_nl = MUX_s_1_2_2((mux_10_nl), (nor_38_nl), FpMul_6U_10U_lor_1_lpi_1_dfm_st_3);
  assign or_38_nl = nor_cse | (~ FpMul_6U_10U_else_2_if_acc_itm_6_1) | FpMul_6U_10U_oelse_1_acc_itm_7_1
      | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp | (~ nor_tmp_1);
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_40, (~ main_stage_v_1), reg_chn_o_rsci_ld_core_psct_cse);
  assign mux_19_nl = MUX_s_1_2_2((mux_18_nl), or_tmp_40, chn_o_rsci_bawt);
  assign mux_20_nl = MUX_s_1_2_2((mux_19_nl), (or_38_nl), or_65_cse);
  assign FpMul_6U_10U_xor_1_nl = (chn_a_rsci_d_mxwt[16]) ^ (chn_b_rsci_d_mxwt[16]);
  assign mux_25_nl = MUX_s_1_2_2(or_tmp_48, (~ nor_tmp_1), FpMul_6U_10U_else_2_if_acc_itm_6_1);
  assign mux_26_nl = MUX_s_1_2_2((mux_25_nl), or_tmp_48, or_68_cse);
  assign mux_27_nl = MUX_s_1_2_2(or_tmp_49, (~ main_stage_v_1), IsNaN_6U_10U_1_land_lpi_1_dfm_3);
  assign mux_28_nl = MUX_s_1_2_2((mux_27_nl), or_tmp_49, IsNaN_6U_10U_land_lpi_1_dfm_st_3);
  assign mux_29_nl = MUX_s_1_2_2((mux_28_nl), (mux_26_nl), or_5_cse);
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_52, nand_6_cse, FpMul_6U_10U_else_2_if_acc_itm_6_1);
  assign mux_31_nl = MUX_s_1_2_2((mux_30_nl), or_tmp_52, or_68_cse);
  assign nor_33_nl = ~(FpMul_6U_10U_lor_1_lpi_1_dfm_st_3 | nand_7_cse);
  assign mux_32_nl = MUX_s_1_2_2((nor_33_nl), main_stage_v_1, IsNaN_6U_10U_land_lpi_1_dfm_st_3);
  assign mux_33_nl = MUX_s_1_2_2((mux_32_nl), (~ (mux_31_nl)), or_5_cse);

  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [9:0] signext_10_1;
    input [0:0] vector;
  begin
    signext_10_1= {{9{vector[0]}}, vector};
  end
  endfunction


  function  [7:0] conv_s2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction


  function  [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function  [7:0] conv_u2s_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [9:0] conv_u2u_1_10 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function  [21:0] conv_u2u_22_22 ;
    input [21:0]  vector ;
  begin
    conv_u2u_22_22 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_mul
// ------------------------------------------------------------------


module HLS_fp17_mul (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;


  // Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_b_rsci_oswt;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;
  wire chn_a_rsci_oswt_unreg_iff;


  // Interconnect Declarations for Component Instantiations 
  FP17_MUL_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_a_rsci_oswt)
    );
  FP17_MUL_chn_b_rsci_unreg chn_b_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_b_rsci_oswt)
    );
  FP17_MUL_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_fp17_mul_core HLS_fp17_mul_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg),
      .chn_a_rsci_oswt_unreg_pff(chn_a_rsci_oswt_unreg_iff)
    );
endmodule



